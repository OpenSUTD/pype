module bannerpart1_7 (
    input wire clk,  // clock
    input wire [7:0] address,  // reset
    output reg [56:0] outdata
  );
  
  (* rom_style = "block" *)
  
  reg [7:0] address_reg;

  /* Combinational Logic */
  always @* begin
    case (address_reg)
        0: outdata = 57'b000000000000000000000000000000000000000000000000000000111;
        1: outdata = 57'b000000000000000000000000000000000000000000000000000000111;
        2: outdata = 57'b000000000000000000000000000000000000000000000000000000111;
        3: outdata = 57'b000000000000000000000000000000000000000000000000111111000;
        4: outdata = 57'b000000000000000000000000000000000000000000000000111111000;
        5: outdata = 57'b000000000000000000000000000000000000000000000000111111000;
        6: outdata = 57'b000000000000000000000000000000000000000000000111000000000;
        7: outdata = 57'b000000000000000000000000000000000000000000000111000000000;
        8: outdata = 57'b000000000000000000000000000000000000000000000111000000000;
        9: outdata = 57'b000000000000000000000000000000000000000111111000000000000;
        10: outdata = 57'b000000000000000000000000000000000000000111111000000000000;
        11: outdata = 57'b000000000000000000000000000000000000000111111000000000000;
        12: outdata = 57'b000000000000000000000000000000000111111000000000000000000;
        13: outdata = 57'b000000000000000000000000000000000111111000000000000000000;
        14: outdata = 57'b000000000000000000000000000000000111111000000000000000000;
        15: outdata = 57'b000000000000000000000000000111111000000000000000000000000;
        16: outdata = 57'b000000000000000000000000000111111000000000000000000000000;
        17: outdata = 57'b000000000000000000000000000111111000000000000000000000000;
        18: outdata = 57'b000000000000000000000000111000000000000000000000000000000;
        19: outdata = 57'b000000000000000000000000111000000000000000000000000000000;
        20: outdata = 57'b000000000000000000000000111000000000000000000000000000000;
        21: outdata = 57'b000000000000000000111111000000000000000000000000000000000;
        22: outdata = 57'b000000000000000000111111000000000000000000000000000000000;
        23: outdata = 57'b000000000000000000111111000000000000000000000000000000000;
        24: outdata = 57'b000000000000111111000000000000000000000000000000000000000;
        25: outdata = 57'b000000000000111111000000000000000000000000000000000000000;
        26: outdata = 57'b000000000000111111000000000000000000000000000000000000000;
        27: outdata = 57'b000000111111000000000000000000000000000000000000000000000;
        28: outdata = 57'b000000111111000000000000000000000000000000000000000000000;
        29: outdata = 57'b000000111111000000000000000000000000000000000000000000000;
        30: outdata = 57'b111111000000000000000000000000000000000000000000000000000;
        31: outdata = 57'b111111000000000000000000000000000000000000000000000000000;
        32: outdata = 57'b111111000000000000000000000000000000000000000000000000000;
        33: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        34: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        35: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        36: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        37: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        38: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        39: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        40: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        41: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        42: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        43: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        44: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        45: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        46: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        47: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        48: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        49: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        50: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        51: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        52: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        53: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        54: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        55: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        56: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        57: outdata = 57'b111000000000000000111111111111000000000000111000000111000;
        58: outdata = 57'b111000000000000000111111111111000000000000111000000111000;
        59: outdata = 57'b111000000000000000111111111111000000000000111000000111000;
        60: outdata = 57'b111000000000000000111111000000111000000000111000000111000;
        61: outdata = 57'b111000000000000000111111000000111000000000111000000111000;
        62: outdata = 57'b111000000000000000111111000000111000000000111000000111000;
        63: outdata = 57'b111000000000000000111111000000111000000000111111111111000;
        64: outdata = 57'b111000000000000000111111000000111000000000111111111111000;
        65: outdata = 57'b111000000000000000111111000000111000000000111111111111000;
        66: outdata = 57'b111000000000000000111111111111000000000000000000111111000;
        67: outdata = 57'b111000000000000000111111111111000000000000000000111111000;
        68: outdata = 57'b111000000000000000111111111111000000000000000000111111000;
        69: outdata = 57'b111000000000000000111111000000000000000000000000111111000;
        70: outdata = 57'b111000000000000000111111000000000000000000000000111111000;
        71: outdata = 57'b111000000000000000111111000000000000000000000000111111000;
        72: outdata = 57'b111000000000000000111111000000000000000000111111111000000;
        73: outdata = 57'b111000000000000000111111000000000000000000111111111000000;
        74: outdata = 57'b111000000000000000111111000000000000000000111111111000000;
        75: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        76: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        77: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        78: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        79: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        80: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        81: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        82: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        83: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        84: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        85: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        86: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        87: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        88: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        89: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        90: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        91: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        92: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        93: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        94: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        95: outdata = 57'b111000000000000000000000000000000000000000000000000000000;
        96: outdata = 57'b000111000000000000000000000000000000000000000000000000000;
        97: outdata = 57'b000111000000000000000000000000000000000000000000000000000;
        98: outdata = 57'b000111000000000000000000000000000000000000000000000000000;
        99: outdata = 57'b000000111111000000000000000000000000000000000000000000000;
        100: outdata = 57'b000000111111000000000000000000000000000000000000000000000;
        101: outdata = 57'b000000111111000000000000000000000000000000000000000000000;
        102: outdata = 57'b000000000000111111000000000000000000000000000000000000000;
        103: outdata = 57'b000000000000111111000000000000000000000000000000000000000;
        104: outdata = 57'b000000000000111111000000000000000000000000000000000000000;
        105: outdata = 57'b000000000000000000111111000000000000000000000000000000000;
        106: outdata = 57'b000000000000000000111111000000000000000000000000000000000;
        107: outdata = 57'b000000000000000000111111000000000000000000000000000000000;
        108: outdata = 57'b000000000000000000000000111000000000000000000000000000000;
        109: outdata = 57'b000000000000000000000000111000000000000000000000000000000;
        110: outdata = 57'b000000000000000000000000111000000000000000000000000000000;
        111: outdata = 57'b000000000000000000000000000111111000000000000000000000000;
        112: outdata = 57'b000000000000000000000000000111111000000000000000000000000;
        113: outdata = 57'b000000000000000000000000000111111000000000000000000000000;
        114: outdata = 57'b000000000000000000000000000000000111111000000000000000000;
        115: outdata = 57'b000000000000000000000000000000000111111000000000000000000;
        116: outdata = 57'b000000000000000000000000000000000111111000000000000000000;
        117: outdata = 57'b000000000000000000000000000000000000000111111000000000000;
        118: outdata = 57'b000000000000000000000000000000000000000111111000000000000;
        119: outdata = 57'b000000000000000000000000000000000000000111111000000000000;
        120: outdata = 57'b000000000000000000000000000000000000000000000111000000000;
        121: outdata = 57'b000000000000000000000000000000000000000000000111000000000;
        122: outdata = 57'b000000000000000000000000000000000000000000000111000000000;
        123: outdata = 57'b000000000000000000000000000000000000000000000000111111000;
        124: outdata = 57'b000000000000000000000000000000000000000000000000111111000;
        125: outdata = 57'b000000000000000000000000000000000000000000000000111111000;
        126: outdata = 57'b000000000000000000000000000000000000000000000000000000111;
        127: outdata = 57'b000000000000000000000000000000000000000000000000000000111;
        128: outdata = 57'b000000000000000000000000000000000000000000000000000000111;


        
        default: outdata = 57'b000000000000000000000000000000000000000000000000000000000000000;
        
        endcase


  end
  
  /* Sequential Logic */
  always @(posedge clk) begin
    address_reg <= address;
  end
  
endmodule
