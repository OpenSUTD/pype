module water (clk, en, address, bitmap);
    input clk;
    input en;
    input wire[5:0] address;
    output reg[589:0] bitmap;
    reg [5:0]address_reg;
    
 always @(posedge clk)
 begin
    if (en)
     address_reg <= address;
 end
 
 always @(address_reg)
 begin
   if(en)
     case(address_reg)
       default: bitmap <= 0;
       6'b000000: bitmap <= 590'b11111100000000000000000000000000000000000000000000000000000000000000000000000000111100000000111111000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000001110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000011110000000011111100000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000111000000000111;
       6'b000001: bitmap <= 590'b11111111100000000000000000011100000000000000011111111100000000000000000000000111111111111111111111111000000000000000000111000000000000000111111111111111111000000000000000000111000000000000000111111111111111110000000000000000001110000000000000001111111110000000000000000000000001111111111111111111111111110000000000000000011110000000000000001111111100000000000000000000000001111111111111111111111100000000000000000011100000000000000011111111111111111100000000000000000011100000000000000111111111111111111000000000000000000111100000000000000111111111000000000000000000000000111111111111111111;
       6'b000010: bitmap <= 590'b11111111111100000000011111111111111111111111100011100011111100000000000000000011111111111111000011111111000000000011111111111111111111111111000111111111111111000000000111111111111111111111111111000111000111111111000000000111111111111111111111111110001111111110000000000000000001111111111111111111111111111110000000001111111111111111111111110001110011111110000000000000000011111111111111100011111111100000000011111111111111111111111111100011111111111111100000000011111111111111111111111111000011100011111111100000000011111111111111111111111111000111111111100000000000000000011111111111111111;
       6'b000011: bitmap <= 590'b00011111111111111111111111111111111100011111111111111111111111111111111111111111111000011000111100111111111111111111111111111111000111111111000111000011111111111111111111111111111111000111111110000111110000111111111111111111111111111110001111111110000111000111111111111111111111111110001110001110001111111111111111111111111111111110001111111111111111111111111111111111111111111100011100001100011111111111111111111111111111100001111111100011100011111111111111111111111111111111100011111111100011111000011111111111111111111111111111000111111111000011100011111111111111111111111111000111000111;
       6'b000100: bitmap <= 590'b00011100000011111111000011100011111111111111100000011100000111111111111000111111111000111111111111000000111111111000111000111111111111110000111111001111000111000111111001111000111111111111110001111111111111000000111111110001110001111111111111110001111110010110001111110001111110001110001111110000001110000001111111100001100001111111111111110000001110000001111111111100011111111100001111111111100000011111111100011100011111111111111100011111100011100011100011111100011100011111111111111000111111111111100000111111111000011000011111111111110100111110001011000011111000111111000111000011111000;
       
       6'b001000: bitmap <= 590'b00000011000000000000000000000000000000000000000000000000000000000000000000000000001111000000001111110000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000011100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000111100000000111111000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000001110000000001;
       6'b001001: bitmap <= 590'b00001111111000000000000000000111000000000000000111111111000000000000000000000001111111111111111111111110000000000000000001110000000000000001111111111111111110000000000000000001110000000000000001111111111111111100000000000000000011100000000000000011111111100000000000000000000000011111111111111111111111111100000000000000000111100000000000000011111111000000000000000000000000011111111111111111111111000000000000000000111000000000000000111111111111111111000000000000000000111000000000000001111111111111111110000000000000000001111000000000000001111111110000000000000000000000001111111111111111;
       6'b001010: bitmap <= 590'b01111111111111000000000111111111111111111111111000111000111111000000000000000000111111111111110000111111110000000000111111111111111111111111110001111111111111110000000001111111111111111111111111110001110001111111110000000001111111111111111111111111100011111111100000000000000000011111111111111111111111111111100000000011111111111111111111111100011100111111100000000000000000111111111111111000111111111000000000111111111111111111111111111000111111111111111000000000111111111111111111111111110000111000111111111000000000111111111111111111111111110001111111111000000000000000000111111111111111;
       6'b001011: bitmap <= 590'b11000111111111111111111111111111111111000111111111111111111111111111111111111111111110000110001111001111111111111111111111111111110001111111110001110000111111111111111111111111111111110001111111100001111100001111111111111111111111111111100011111111100001110001111111111111111111111111100011100011100011111111111111111111111111111111100011111111111111111111111111111111111111111111000111000011000111111111111111111111111111111000011111111000111000111111111111111111111111111111111000111111111000111110000111111111111111111111111111110001111111110000111000111111111111111111111111110001110001;
       6'b001100: bitmap <= 590'b11000111000000111111110000111000111111111111111000000111000001111111111110001111111110001111111111110000001111111110001110001111111111111100001111110011110001110001111110011110001111111111111100011111111111110000001111111100011100011111111111111100011111100101100011111100011111100011100011111100000011100000011111111000011000011111111111111100000011100000011111111111000111111111000011111111111000000111111111000111000111111111111111000111111000111000111000111111000111000111111111111110001111111111111000001111111110000110000111111111111101001111100010110000111110001111110001110000111110;

       6'b010000: bitmap <= 590'b11110000000000000000000000000000000000000000000000000000000000000000000000000011110000000011111100000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000001111000000001111110000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000;
       6'b010001: bitmap <= 590'b11111110000000000000000001110000000000000001111111110000000000000000000000011111111111111111111111100000000000000000011100000000000000011111111111111111100000000000000000011100000000000000011111111111111111000000000000000000111000000000000000111111111000000000000000000000000111111111111111111111111111000000000000000001111000000000000000111111110000000000000000000000000111111111111111111111110000000000000000001110000000000000001111111111111111110000000000000000001110000000000000011111111111111111100000000000000000011110000000000000011111111100000000000000000000000011111111111111110000;
       6'b010010: bitmap <= 590'b11111111110000000001111111111111111111111110001110001111110000000000000000001111111111111100001111111100000000001111111111111111111111111100011111111111111100000000011111111111111111111111111100011100011111111100000000011111111111111111111111111000111111111000000000000000000111111111111111111111111111111000000000111111111111111111111111000111001111111000000000000000001111111111111110001111111110000000001111111111111111111111111110001111111111111110000000001111111111111111111111111100001110001111111110000000001111111111111111111111111100011111111110000000000000000001111111111111111100;
       6'b010011: bitmap <= 590'b01111111111111111111111111111111110001111111111111111111111111111111111111111111100001100011110011111111111111111111111111111100011111111100011100001111111111111111111111111111111100011111111000011111000011111111111111111111111111111000111111111000011100011111111111111111111111111000111000111000111111111111111111111111111111111000111111111111111111111111111111111111111111110001110000110001111111111111111111111111111110000111111110001110001111111111111111111111111111111110001111111110001111100001111111111111111111111111111100011111111100001110001111111111111111111111111100011100011111;
       6'b010100: bitmap <= 590'b01110000001111111100001110001111111111111110000001110000011111111111100011111111100011111111111100000011111111100011100011111111111111000011111100111100011100011111100111100011111111111111000111111111111100000011111111000111000111111111111111000111111001011000111111000111111000111000111111000000111000000111111110000110000111111111111111000000111000000111111111110001111111110000111111111110000001111111110001110001111111111111110001111110001110001110001111110001110001111111111111100011111111111110000011111111100001100001111111111111010011111000101100001111100011111100011100001111100011;
     endcase
 end
  
endmodule
