module selector_base_36 (
    input wire clk,  // clock
    input wire[6:0] address,
    output reg [58:0] outdata
  );
  
  (* rom_style = "block" *)
  
  reg [6:0] address_reg;

  /* Combinational Logic */
  always @* begin
    case(address)
      0: outdata = 59'b00000000000000000000000000111111100000000000000000000000000;
      1: outdata = 59'b00000000000000000000000011111111111000000000000000000000000;
      2: outdata = 59'b00000000000000000000001111100000111110000000000000000000000;
      3: outdata = 59'b00000000000000000000011110000000001111000000000000000000000;
      4: outdata = 59'b00000000000000000001111000000000000011110000000000000000000;
      5: outdata = 59'b00000000000000000011110000000000000001111000000000000000000;
      6: outdata = 59'b00000000000000001111000000000000000000011110000000000000000;
      7: outdata = 59'b00000000000000111100000000000000000000000111100000000000000;
      8: outdata = 59'b00000000000001111000000000000000000000000011110000000000000;
      9: outdata = 59'b00000000000111100000000000000000000000000000111100000000000;
      10: outdata = 59'b00000000011110000000000000000000000000000000001111000000000;
      11: outdata = 59'b00000000111000000000000000000000000000000000000011100000000;
      12: outdata = 59'b00000011110000000000000000000000000000000000000001111000000;
      13: outdata = 59'b00000111000000000000000000000000000000000000000000011100000;
      14: outdata = 59'b00011100000000000000000000000000000000000000000000000111000;
      15: outdata = 59'b01111000000000000000000000000000000000000000000000000011110;
      16: outdata = 59'b01100000000000000000000000000000000000000000000000000000110;
      17: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      18: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      19: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      20: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      21: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      22: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      23: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      24: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      25: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      26: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      27: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      28: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      29: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      30: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      31: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      32: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      33: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      34: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      35: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      36: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      37: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      38: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      39: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      40: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      41: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      42: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      43: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      44: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      45: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      46: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      47: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      48: outdata = 59'b11000000000000000000000000000000000000000000000000000000011;
      49: outdata = 59'b01100000000000000000000000000000000000000000000000000000110;
      50: outdata = 59'b01111000000000000000000000000000000000000000000000000011110;
      51: outdata = 59'b00011100000000000000000000000000000000000000000000000111000;
      52: outdata = 59'b00000111000000000000000000000000000000000000000000011100000;
      53: outdata = 59'b00000011110000000000000000000000000000000000000001111000000;
      54: outdata = 59'b00000000111000000000000000000000000000000000000011100000000;
      55: outdata = 59'b00000000011110000000000000000000000000000000001111000000000;
      56: outdata = 59'b00000000000111100000000000000000000000000000111100000000000;
      57: outdata = 59'b00000000000001111000000000000000000000000011110000000000000;
      58: outdata = 59'b00000000000000111100000000000000000000000111100000000000000;
      59: outdata = 59'b00000000000000001111000000000000000000011110000000000000000;
      60: outdata = 59'b00000000000000000011110000000000000001111000000000000000000;
      61: outdata = 59'b00000000000000000001111000000000000011110000000000000000000;
      62: outdata = 59'b00000000000000000000011110000000001111000000000000000000000;
      63: outdata = 59'b00000000000000000000001111100000111110000000000000000000000;
      64: outdata = 59'b00000000000000000000000011111111111000000000000000000000000;
      65: outdata = 59'b00000000000000000000000000111111100000000000000000000000000;    
    endcase
  end
  
  /* Sequential Logic */
  always @(posedge clk) begin
    address_reg <= address;    
  end
  
endmodule