module tile_library (
    input wire clk,  // clock
    input wire[5:0] data,
    input wire[5:0] address,
    output reg[50:0] bitmap
  );
  
  (* rom_style = "block" *)

  reg[5:0] data_reg;  
  reg[5:0] address_reg;
  
  always @(posedge clk) begin
    address_reg <= address;
    data_reg <= data;
    
  end

  /* Combinational Logic */
  always @* begin
      case({data_reg,address_reg})
        default: bitmap = 0;
        12'b000000000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b000000000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b000000000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b000000000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b000000000100: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b000000000101: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b000000000110: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b000000000111: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b000000001000: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b000000001001: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b000000001010: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b000000001011: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b000000001100: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b000000001101: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b000000001110: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b000000001111: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b000000010000: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b000000010001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b000000010010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b000000010011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b000000010100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b000000010101: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b000000010110: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b000000010111: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b000000011000: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b000000011001: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b000000011010: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b000000011011: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b000000011100: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b000000011101: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b000000011110: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b000000011111: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b000000100000: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b000000100001: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b000000100010: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b000000100011: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b000000100100: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b000000100101: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b000000100110: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b000000100111: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b000000101000: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b000000101001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b000000101010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b000000101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b000000101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b000000101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b000000101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b000000101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b000000110000: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b000000110001: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b000000110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b000000110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b000000110100: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b000000110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b000000110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b000000110111: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b000000111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b000000111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b000000111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b000000111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        
        
        12'b000001000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b000001000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b000001000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b000001000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b000001000100: bitmap = 51'b000000000000000000011111111111111000000000000000000;
        12'b000001000101: bitmap = 51'b000000000000000000001111111111111110000000000000000;
        12'b000001000110: bitmap = 51'b000000000000000000001111111111111111100000000000000;
        12'b000001000111: bitmap = 51'b000000000000000000000111111111111111110000000000000;
        12'b000001001000: bitmap = 51'b000000000000000000000111111111111111111100000000000;
        12'b000001001001: bitmap = 51'b000000000000000000000011111111111111111111000000000;
        12'b000001001010: bitmap = 51'b000000000000000000000011111111111111111111100000000;
        12'b000001001011: bitmap = 51'b000000100000000000000001111111111111111111111000000;
        12'b000001001100: bitmap = 51'b000011110000000000000000111111111111111111111110000;
        12'b000001001101: bitmap = 51'b000111110000000000000000111111111111111111111111000;
        12'b000001001110: bitmap = 51'b011111111000000000000000011111111111111111111111110;
        12'b000001001111: bitmap = 51'b111111111000000000000000011111111111111111111111111;
        12'b000001010000: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b000001010001: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b000001010010: bitmap = 51'b111111111110000000000000000111111111111111111111111;
        12'b000001010011: bitmap = 51'b111111111111000000000000000011111111111111111111111;
        12'b000001010100: bitmap = 51'b111111111111000000000000000011111111111111111111111;
        12'b000001010101: bitmap = 51'b111111111111100000000000000001111111111111111111111;
        12'b000001010110: bitmap = 51'b111111111111100000000000000001111111111111111111111;
        12'b000001010111: bitmap = 51'b111111111111110000000000000000111111111111111111111;
        12'b000001011000: bitmap = 51'b111111111111110000000000000000111111111111111111111;
        12'b000001011001: bitmap = 51'b111111111111111000000000000000011111111111111111111;
        12'b000001011010: bitmap = 51'b111111111111111100000000000000011111111111111111111;
        12'b000001011011: bitmap = 51'b111111111111111100000000000000001111111111111111111;
        12'b000001011100: bitmap = 51'b111111111111111110000000000000000111111111111111111;
        12'b000001011101: bitmap = 51'b111111111111111110000000000000000111111111111111111;
        12'b000001011110: bitmap = 51'b111111111111111111000000000000000011111111111111111;
        12'b000001011111: bitmap = 51'b111111111111111111000000000000000011111111111111111;
        12'b000001100000: bitmap = 51'b111111111111111111100000000000000001111111111111111;
        12'b000001100001: bitmap = 51'b111111111111111111100000000000000001111111111111111;
        12'b000001100010: bitmap = 51'b111111111111111111110000000000000000111111111111111;
        12'b000001100011: bitmap = 51'b111111111111111111111000000000000000011111111111111;
        12'b000001100100: bitmap = 51'b111111111111111111111000000000000000011111111111111;
        12'b000001100101: bitmap = 51'b111111111111111111111100000000000000001111111111111;
        12'b000001100110: bitmap = 51'b111111111111111111111100000000000000001111111111111;
        12'b000001100111: bitmap = 51'b111111111111111111111110000000000000000111111111111;
        12'b000001101000: bitmap = 51'b111111111111111111111110000000000000000111111111111;
        12'b000001101001: bitmap = 51'b111111111111111111111111000000000000000011111111111;
        12'b000001101010: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b000001101011: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b000001101100: bitmap = 51'b111111111111111111111111110000000000000000111111111;
        12'b000001101101: bitmap = 51'b011111111111111111111111110000000000000000111111110;
        12'b000001101110: bitmap = 51'b000111111111111111111111111000000000000000011111000;
        12'b000001101111: bitmap = 51'b000011111111111111111111111000000000000000011110000;
        12'b000001110000: bitmap = 51'b000000111111111111111111111100000000000000001000000;
        12'b000001110001: bitmap = 51'b000000001111111111111111111110000000000000000000000;
        12'b000001110010: bitmap = 51'b000000000111111111111111111110000000000000000000000;
        12'b000001110011: bitmap = 51'b000000000001111111111111111111000000000000000000000;
        12'b000001110100: bitmap = 51'b000000000000011111111111111111000000000000000000000;
        12'b000001110101: bitmap = 51'b000000000000001111111111111111100000000000000000000;
        12'b000001110110: bitmap = 51'b000000000000000011111111111111100000000000000000000;
        12'b000001110111: bitmap = 51'b000000000000000000111111111111110000000000000000000;
        12'b000001111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b000001111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b000001111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b000001111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        
        //shape 1
        12'b001000000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b001000000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b001000000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b001000000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b001000000100: bitmap = 51'b000000000000000000111111111111110000000000000000000;
        12'b001000000101: bitmap = 51'b000000000000000011111111111111100000000000000000000;
        12'b001000000110: bitmap = 51'b000000000000001111111111111111100000000000000000000;
        12'b001000000111: bitmap = 51'b000000000000011111111111111111000000000000000000000;
        12'b001000001000: bitmap = 51'b000000000001111111111111111111000000000000000000000;
        12'b001000001001: bitmap = 51'b000000000111111111111111111110000000000000000000000;
        12'b001000001010: bitmap = 51'b000000001111111111111111111110000000000000000000000;
        12'b001000001011: bitmap = 51'b000000111111111111111111111100000000000000001000000;
        12'b001000001100: bitmap = 51'b000011111111111111111111111000000000000000011110000;
        12'b001000001101: bitmap = 51'b000111111111111111111111111000000000000000011111000;
        12'b001000001110: bitmap = 51'b011111111111111111111111110000000000000000111111110;
        12'b001000001111: bitmap = 51'b111111111111111111111111110000000000000000111111111;
        12'b001000010000: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b001000010001: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b001000010010: bitmap = 51'b111111111111111111111111000000000000000011111111111;
        12'b001000010011: bitmap = 51'b111111111111111111111110000000000000000111111111111;
        12'b001000010100: bitmap = 51'b111111111111111111111110000000000000000111111111111;
        12'b001000010101: bitmap = 51'b111111111111111111111100000000000000001111111111111;
        12'b001000010110: bitmap = 51'b111111111111111111110000000000000000001111111111111;
        12'b001000010111: bitmap = 51'b000000000000000000000000000000000000011111111111111;
        12'b001000011000: bitmap = 51'b000000000000000000000000000000000000011111111111111;
        12'b001000011001: bitmap = 51'b000000000000000000000000000000000000111111111111111;
        12'b001000011010: bitmap = 51'b000000000000000000000000000000000001111111111111111;
        12'b001000011011: bitmap = 51'b000000000000000000000000000000000001111111111111111;
        12'b001000011100: bitmap = 51'b000000000000000000000000000000000011111111111111111;
        12'b001000011101: bitmap = 51'b000000000000000000000000000000000011111111111111111;
        12'b001000011110: bitmap = 51'b000000000000000000000000000000000111111111111111111;
        12'b001000011111: bitmap = 51'b000000000000000000000000000000000111111111111111111;
        12'b001000100000: bitmap = 51'b000000000000000000000000000000001111111111111111111;
        12'b001000100001: bitmap = 51'b000000000000000000000000000000011111111111111111111;
        12'b001000100010: bitmap = 51'b000000000000000000000000000000111111111111111111111;
        12'b001000100011: bitmap = 51'b000000000000000000000000000011111111111111111111111;
        12'b001000100100: bitmap = 51'b000000000000000000000000001111111111111111111111111;
        12'b001000100101: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b001000100110: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b001000100111: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b001000101000: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b001000101001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b001000101010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b001000101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b001000101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b001000101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b001000101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b001000101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b001000110000: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b001000110001: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b001000110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b001000110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b001000110100: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b001000110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b001000110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b001000110111: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b001000111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b001000111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b001000111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b001000111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;




        
        12'b001001000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b001001000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b001001000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b001001000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b001001000100: bitmap = 51'b000000000000000000011111111111111000000000000000000;
        12'b001001000101: bitmap = 51'b000000000000000000001111111111111110000000000000000;
        12'b001001000110: bitmap = 51'b000000000000000000001111111111111111100000000000000;
        12'b001001000111: bitmap = 51'b000000000000000000000111111111111111110000000000000;
        12'b001001001000: bitmap = 51'b000000000000000000000111111111111111111100000000000;
        12'b001001001001: bitmap = 51'b000000000000000000000011111111111111111111000000000;
        12'b001001001010: bitmap = 51'b000000000000000000000011111111111111111111100000000;
        12'b001001001011: bitmap = 51'b000000100000000000000001111111111111111111111000000;
        12'b001001001100: bitmap = 51'b000011110000000000000000111111111111111111111110000;
        12'b001001001101: bitmap = 51'b000111110000000000000000111111111111111111111111000;
        12'b001001001110: bitmap = 51'b011111111000000000000000011111111111111111111111110;
        12'b001001001111: bitmap = 51'b111111111000000000000000011111111111111111111111111;
        12'b001001010000: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b001001010001: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b001001010010: bitmap = 51'b111111111110000000000000000111111111111111111111111;
        12'b001001010011: bitmap = 51'b111111111111000000000000000011111111111111111111111;
        12'b001001010100: bitmap = 51'b111111111111000000000000000011111111111111111111111;
        12'b001001010101: bitmap = 51'b111111111111100000000000000001111111111111111111111;
        12'b001001010110: bitmap = 51'b111111111111100000000000000000011111111111111111111;
        12'b001001010111: bitmap = 51'b111111111111110000000000000000000000000000000000000;
        12'b001001011000: bitmap = 51'b111111111111110000000000000000000000000000000000000;
        12'b001001011001: bitmap = 51'b111111111111111000000000000000000000000000000000000;
        12'b001001011010: bitmap = 51'b111111111111111100000000000000000000000000000000000;
        12'b001001011011: bitmap = 51'b111111111111111100000000000000000000000000000000000;
        12'b001001011100: bitmap = 51'b111111111111111110000000000000000000000000000000000;
        12'b001001011101: bitmap = 51'b111111111111111110000000000000000000000000000000000;
        12'b001001011110: bitmap = 51'b111111111111111111000000000000000000000000000000000;
        12'b001001011111: bitmap = 51'b111111111111111111000000000000000000000000000000000;
        12'b001001100000: bitmap = 51'b111111111111111111100000000000000000000000000000000;
        12'b001001100001: bitmap = 51'b111111111111111111110000000000000000000000000000000;
        12'b001001100010: bitmap = 51'b111111111111111111111000000000000000000000000000000;
        12'b001001100011: bitmap = 51'b111111111111111111111110000000000000000000000000000;
        12'b001001100100: bitmap = 51'b111111111111111111111111100000000000000000000000000;
        12'b001001100101: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b001001100110: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b001001100111: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b001001101000: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b001001101001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b001001101010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b001001101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b001001101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b001001101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b001001101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b001001101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b001001110000: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b001001110001: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b001001110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b001001110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b001001110100: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b001001110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b001001110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b001001110111: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b001001111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b001001111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b001001111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b001001111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;


        
        12'b001010000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b001010000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b001010000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b001010000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b001010000100: bitmap = 51'b000000000000000000011111111111100000000000000000000;
        12'b001010000101: bitmap = 51'b000000000000000011111111111111100000000000000000000;
        12'b001010000110: bitmap = 51'b000000000000001111111111111111000000000000000000000;
        12'b001010000111: bitmap = 51'b000000000000011111111111111111000000000000000000000;
        12'b001010001000: bitmap = 51'b000000000001111111111111111110000000000000000000000;
        12'b001010001001: bitmap = 51'b000000000111111111111111111110000000000000000000000;
        12'b001010001010: bitmap = 51'b000000001111111111111111111100000000000000000000000;
        12'b001010001011: bitmap = 51'b000000111111111111111111111100000000000000001000000;
        12'b001010001100: bitmap = 51'b000011111111111111111111111000000000000000001110000;
        12'b001010001101: bitmap = 51'b000111111111111111111111110000000000000000011111000;
        12'b001010001110: bitmap = 51'b011111111111111111111111110000000000000000111111110;
        12'b001010001111: bitmap = 51'b111111111111111111111111100000000000000000111111111;
        12'b001010010000: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b001010010001: bitmap = 51'b111111111111111111111111000000000000000001111111111;
        12'b001010010010: bitmap = 51'b111111111111111111111111000000000000000011111111111;
        12'b001010010011: bitmap = 51'b111111111111111111111110000000000000000111111111111;
        12'b001010010100: bitmap = 51'b111111111111111111111110000000000000000111111111111;
        12'b001010010101: bitmap = 51'b111111111111111111111100000000000000001111111111111;
        12'b001010010110: bitmap = 51'b111111111111111111111000000000000000001111111111111;
        12'b001010010111: bitmap = 51'b111111111111111111111000000000000000011111111111111;
        12'b001010011000: bitmap = 51'b111111111111111111110000000000000000011111111111111;
        12'b001010011001: bitmap = 51'b111111111111111111110000000000000000111111111111111;
        12'b001010011010: bitmap = 51'b111111111111111111100000000000000001111111111111111;
        12'b001010011011: bitmap = 51'b111111111111111111100000000000000001111111111111111;
        12'b001010011100: bitmap = 51'b111111111111111111100000000000000001111111111111111;
        12'b001010011101: bitmap = 51'b111111111111111111100000000000000011111111111111111;
        12'b001010011110: bitmap = 51'b111111111111111111100000000000000011111111111111111;
        12'b001010011111: bitmap = 51'b111111111111111111100000000000000001111111111111111;
        12'b001010100000: bitmap = 51'b111111111111111111100000000000000001111111111111111;
        12'b001010100001: bitmap = 51'b111111111111111111110000000000000001111111111111111;
        12'b001010100010: bitmap = 51'b111111111111111111110000000000000000111111111111111;
        12'b001010100011: bitmap = 51'b111111111111111111111000000000000000011111111111111;
        12'b001010100100: bitmap = 51'b111111111111111111111000000000000000011111111111111;
        12'b001010100101: bitmap = 51'b111111111111111111111100000000000000001111111111111;
        12'b001010100110: bitmap = 51'b111111111111111111111110000000000000001111111111111;
        12'b001010100111: bitmap = 51'b111111111111111111111110000000000000000111111111111;
        12'b001010101000: bitmap = 51'b111111111111111111111111000000000000000111111111111;
        12'b001010101001: bitmap = 51'b111111111111111111111111000000000000000011111111111;
        12'b001010101010: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b001010101011: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b001010101100: bitmap = 51'b111111111111111111111111110000000000000000111111111;
        12'b001010101101: bitmap = 51'b011111111111111111111111110000000000000000111111110;
        12'b001010101110: bitmap = 51'b000111111111111111111111111000000000000000011111000;
        12'b001010101111: bitmap = 51'b000011111111111111111111111100000000000000011110000;
        12'b001010110000: bitmap = 51'b000000111111111111111111111100000000000000001000000;
        12'b001010110001: bitmap = 51'b000000001111111111111111111110000000000000000000000;
        12'b001010110010: bitmap = 51'b000000000111111111111111111110000000000000000000000;
        12'b001010110011: bitmap = 51'b000000000001111111111111111111000000000000000000000;
        12'b001010110100: bitmap = 51'b000000000000011111111111111111000000000000000000000;
        12'b001010110101: bitmap = 51'b000000000000001111111111111111100000000000000000000;
        12'b001010110110: bitmap = 51'b000000000000000011111111111111100000000000000000000;
        12'b001010110111: bitmap = 51'b000000000000000000111111111111110000000000000000000;
        12'b001010111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b001010111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b001010111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b001010111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        
        
        12'b001011000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b001011000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b001011000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b001011000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b001011000100: bitmap = 51'b000000000000000000001111111111110000000000000000000;
        12'b001011000101: bitmap = 51'b000000000000000000001111111111111110000000000000000;
        12'b001011000110: bitmap = 51'b000000000000000000000111111111111111100000000000000;
        12'b001011000111: bitmap = 51'b000000000000000000000111111111111111110000000000000;
        12'b001011001000: bitmap = 51'b000000000000000000000011111111111111111100000000000;
        12'b001011001001: bitmap = 51'b000000000000000000000011111111111111111111000000000;
        12'b001011001010: bitmap = 51'b000000000000000000000001111111111111111111100000000;
        12'b001011001011: bitmap = 51'b000000100000000000000001111111111111111111111000000;
        12'b001011001100: bitmap = 51'b000011100000000000000000111111111111111111111110000;
        12'b001011001101: bitmap = 51'b000111110000000000000000011111111111111111111111000;
        12'b001011001110: bitmap = 51'b011111111000000000000000011111111111111111111111110;
        12'b001011001111: bitmap = 51'b111111111000000000000000001111111111111111111111111;
        12'b001011010000: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b001011010001: bitmap = 51'b111111111100000000000000000111111111111111111111111;
        12'b001011010010: bitmap = 51'b111111111110000000000000000111111111111111111111111;
        12'b001011010011: bitmap = 51'b111111111111000000000000000011111111111111111111111;
        12'b001011010100: bitmap = 51'b111111111111000000000000000011111111111111111111111;
        12'b001011010101: bitmap = 51'b111111111111100000000000000001111111111111111111111;
        12'b001011010110: bitmap = 51'b111111111111100000000000000000111111111111111111111;
        12'b001011010111: bitmap = 51'b111111111111110000000000000000111111111111111111111;
        12'b001011011000: bitmap = 51'b111111111111110000000000000000011111111111111111111;
        12'b001011011001: bitmap = 51'b111111111111111000000000000000011111111111111111111;
        12'b001011011010: bitmap = 51'b111111111111111100000000000000001111111111111111111;
        12'b001011011011: bitmap = 51'b111111111111111100000000000000001111111111111111111;
        12'b001011011100: bitmap = 51'b111111111111111100000000000000001111111111111111111;
        12'b001011011101: bitmap = 51'b111111111111111110000000000000001111111111111111111;
        12'b001011011110: bitmap = 51'b111111111111111110000000000000001111111111111111111;
        12'b001011011111: bitmap = 51'b111111111111111100000000000000001111111111111111111;
        12'b001011100000: bitmap = 51'b111111111111111100000000000000001111111111111111111;
        12'b001011100001: bitmap = 51'b111111111111111100000000000000011111111111111111111;
        12'b001011100010: bitmap = 51'b111111111111111000000000000000011111111111111111111;
        12'b001011100011: bitmap = 51'b111111111111110000000000000000111111111111111111111;
        12'b001011100100: bitmap = 51'b111111111111110000000000000000111111111111111111111;
        12'b001011100101: bitmap = 51'b111111111111100000000000000001111111111111111111111;
        12'b001011100110: bitmap = 51'b111111111111100000000000000011111111111111111111111;
        12'b001011100111: bitmap = 51'b111111111111000000000000000011111111111111111111111;
        12'b001011101000: bitmap = 51'b111111111111000000000000000111111111111111111111111;
        12'b001011101001: bitmap = 51'b111111111110000000000000000111111111111111111111111;
        12'b001011101010: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b001011101011: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b001011101100: bitmap = 51'b111111111000000000000000011111111111111111111111111;
        12'b001011101101: bitmap = 51'b011111111000000000000000011111111111111111111111110;
        12'b001011101110: bitmap = 51'b000111110000000000000000111111111111111111111111000;
        12'b001011101111: bitmap = 51'b000011110000000000000001111111111111111111111110000;
        12'b001011110000: bitmap = 51'b000000100000000000000001111111111111111111111000000;
        12'b001011110001: bitmap = 51'b000000000000000000000011111111111111111111100000000;
        12'b001011110010: bitmap = 51'b000000000000000000000011111111111111111111000000000;
        12'b001011110011: bitmap = 51'b000000000000000000000111111111111111111100000000000;
        12'b001011110100: bitmap = 51'b000000000000000000000111111111111111110000000000000;
        12'b001011110101: bitmap = 51'b000000000000000000001111111111111111100000000000000;
        12'b001011110110: bitmap = 51'b000000000000000000001111111111111110000000000000000;
        12'b001011110111: bitmap = 51'b000000000000000000011111111111111000000000000000000;
        12'b001011111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b001011111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b001011111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b001011111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;

       //shape 2
        12'b010000000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b010000000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b010000000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b010000000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b010000000100: bitmap = 51'b000000000000000000011111111111110000000000000000000;
        12'b010000000101: bitmap = 51'b000000000000000000001111111111111110000000000000000;
        12'b010000000110: bitmap = 51'b000000000000000000001111111111111111100000000000000;
        12'b010000000111: bitmap = 51'b000000000000000000000111111111111111110000000000000;
        12'b010000001000: bitmap = 51'b000000000000000000000111111111111111111100000000000;
        12'b010000001001: bitmap = 51'b000000000000000000000011111111111111111111000000000;
        12'b010000001010: bitmap = 51'b000000000000000000000011111111111111111111100000000;
        12'b010000001011: bitmap = 51'b000000100000000000000001111111111111111111111000000;
        12'b010000001100: bitmap = 51'b000011110000000000000001111111111111111111111110000;
        12'b010000001101: bitmap = 51'b000111110000000000000000111111111111111111111111000;
        12'b010000001110: bitmap = 51'b011111111000000000000000011111111111111111111111110;
        12'b010000001111: bitmap = 51'b111111111000000000000000011111111111111111111111111;
        12'b010000010000: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b010000010001: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b010000010010: bitmap = 51'b111111111110000000000000000111111111111111111111111;
        12'b010000010011: bitmap = 51'b111111111111000000000000000111111111111111111111111;
        12'b010000010100: bitmap = 51'b111111111111000000000000000011111111111111111111111;
        12'b010000010101: bitmap = 51'b111111111111100000000000000011111111111111111111111;
        12'b010000010110: bitmap = 51'b111111111111100000000000000001111111111111111111111;
        12'b010000010111: bitmap = 51'b000000000000000000000000000000111111111111111111111;
        12'b010000011000: bitmap = 51'b000000000000000000000000000000111111111111111111111;
        12'b010000011001: bitmap = 51'b000000000000000000000000000000011111111111111111111;
        12'b010000011010: bitmap = 51'b000000000000000000000000000000011111111111111111111;
        12'b010000011011: bitmap = 51'b000000000000000000000000000000001111111111111111111;
        12'b010000011100: bitmap = 51'b000000000000000000000000000000001111111111111111111;
        12'b010000011101: bitmap = 51'b000000000000000000000000000000001111111111111111111;
        12'b010000011110: bitmap = 51'b000000000000000000000000000000001111111111111111111;
        12'b010000011111: bitmap = 51'b000000000000000000000000000000001111111111111111111;
        12'b010000100000: bitmap = 51'b000000000000000000000000000000001111111111111111111;
        12'b010000100001: bitmap = 51'b000000000000000000000000000000011111111111111111111;
        12'b010000100010: bitmap = 51'b000000000000000000000000000000011111111111111111111;
        12'b010000100011: bitmap = 51'b000000000000000000000000000000111111111111111111111;
        12'b010000100100: bitmap = 51'b000000000000000000000000000000111111111111111111111;
        12'b010000100101: bitmap = 51'b111111111111110000000000000001111111111111111111111;
        12'b010000100110: bitmap = 51'b111111111111100000000000000001111111111111111111111;
        12'b010000100111: bitmap = 51'b111111111111100000000000000011111111111111111111111;
        12'b010000101000: bitmap = 51'b111111111111000000000000000011111111111111111111111;
        12'b010000101001: bitmap = 51'b111111111110000000000000000111111111111111111111111;
        12'b010000101010: bitmap = 51'b111111111110000000000000001111111111111111111111111;
        12'b010000101011: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b010000101100: bitmap = 51'b111111111100000000000000011111111111111111111111111;
        12'b010000101101: bitmap = 51'b011111111000000000000000011111111111111111111111110;
        12'b010000101110: bitmap = 51'b000111111000000000000000111111111111111111111111000;
        12'b010000101111: bitmap = 51'b000011110000000000000000111111111111111111111110000;
        12'b010000110000: bitmap = 51'b000000110000000000000001111111111111111111111000000;
        12'b010000110001: bitmap = 51'b000000000000000000000011111111111111111111100000000;
        12'b010000110010: bitmap = 51'b000000000000000000000011111111111111111111000000000;
        12'b010000110011: bitmap = 51'b000000000000000000000111111111111111111100000000000;
        12'b010000110100: bitmap = 51'b000000000000000000000111111111111111110000000000000;
        12'b010000110101: bitmap = 51'b000000000000000000001111111111111111100000000000000;
        12'b010000110110: bitmap = 51'b000000000000000000001111111111111110000000000000000;
        12'b010000110111: bitmap = 51'b000000000000000000011111111111110000000000000000000;
        12'b010000111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b010000111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b010000111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b010000111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;

        
        12'b010001000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b010001000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b010001000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b010001000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b010001000100: bitmap = 51'b000000000000000000011111111111110000000000000000000;
        12'b010001000101: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b010001000110: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b010001000111: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b010001001000: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b010001001001: bitmap = 51'b000000000000000000000011111110000000000000000000000;
        12'b010001001010: bitmap = 51'b000000000000000000000011111110000000000000000000000;
        12'b010001001011: bitmap = 51'b000000100000000000000001111100000000000000001000000;
        12'b010001001100: bitmap = 51'b000011110000000000000001111100000000000000011110000;
        12'b010001001101: bitmap = 51'b000111110000000000000000111000000000000000011111000;
        12'b010001001110: bitmap = 51'b011111111000000000000000010000000000000000111111110;
        12'b010001001111: bitmap = 51'b111111111000000000000000010000000000000000111111111;
        12'b010001010000: bitmap = 51'b111111111100000000000000000000000000000001111111111;
        12'b010001010001: bitmap = 51'b111111111100000000000000000000000000000001111111111;
        12'b010001010010: bitmap = 51'b111111111110000000000000000000000000000011111111111;
        12'b010001010011: bitmap = 51'b111111111110000000000000000000000000000011111111111;
        12'b010001010100: bitmap = 51'b111111111111000000000000000000000000000111111111111;
        12'b010001010101: bitmap = 51'b111111111111100000000000000000000000001111111111111;
        12'b010001010110: bitmap = 51'b111111111111100000000000000000000000001111111111111;
        12'b010001010111: bitmap = 51'b000000000000000000000000000000000000011111111111111;
        12'b010001011000: bitmap = 51'b000000000000000000000000000000000000011111111111111;
        12'b010001011001: bitmap = 51'b000000000000000000000000000000000000111111111111111;
        12'b010001011010: bitmap = 51'b000000000000000000000000000000000000111111111111111;
        12'b010001011011: bitmap = 51'b000000000000000000000000000000000001111111111111111;
        12'b010001011100: bitmap = 51'b000000000000000000000000000000000001111111111111111;
        12'b010001011101: bitmap = 51'b000000000000000000000000000000000011111111111111111;
        12'b010001011110: bitmap = 51'b000000000000000000000000000000000011111111111111111;
        12'b010001011111: bitmap = 51'b000000000000000000000000000000000111111111111111111;
        12'b010001100000: bitmap = 51'b000000000000000000000000000000001111111111111111111;
        12'b010001100001: bitmap = 51'b000000000000000000000000000000011111111111111111111;
        12'b010001100010: bitmap = 51'b000000000000000000000000000000111111111111111111111;
        12'b010001100011: bitmap = 51'b000000000000000000000000000011111111111111111111111;
        12'b010001100100: bitmap = 51'b000000000000000000000000001111111111111111111111111;
        12'b010001100101: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b010001100110: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b010001100111: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b010001101000: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b010001101001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b010001101010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b010001101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b010001101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b010001101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b010001101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b010001101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b010001110000: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b010001110001: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b010001110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b010001110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b010001110100: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b010001110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b010001110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b010001110111: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b010001111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b010001111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b010001111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b010001111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;

        
        12'b010010000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b010010000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b010010000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b010010000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b010010000100: bitmap = 51'b000000000000000000011111111111110000000000000000000;
        12'b010010000101: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b010010000110: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b010010000111: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b010010001000: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b010010001001: bitmap = 51'b000000000000000000000011111110000000000000000000000;
        12'b010010001010: bitmap = 51'b000000000000000000000011111110000000000000000000000;
        12'b010010001011: bitmap = 51'b000000100000000000000001111100000000000000001000000;
        12'b010010001100: bitmap = 51'b000011110000000000000001111100000000000000011110000;
        12'b010010001101: bitmap = 51'b000111110000000000000000111000000000000000011111000;
        12'b010010001110: bitmap = 51'b011111111000000000000000010000000000000000111111110;
        12'b010010001111: bitmap = 51'b111111111000000000000000010000000000000000111111111;
        12'b010010010000: bitmap = 51'b111111111100000000000000000000000000000001111111111;
        12'b010010010001: bitmap = 51'b111111111100000000000000000000000000000001111111111;
        12'b010010010010: bitmap = 51'b111111111110000000000000000000000000000011111111111;
        12'b010010010011: bitmap = 51'b111111111110000000000000000000000000000011111111111;
        12'b010010010100: bitmap = 51'b111111111111000000000000000000000000000111111111111;
        12'b010010010101: bitmap = 51'b111111111111100000000000000000000000001111111111111;
        12'b010010010110: bitmap = 51'b111111111111100000000000000000000000001111111111111;
        12'b010010010111: bitmap = 51'b111111111111110000000000000000000000000000000000000;
        12'b010010011000: bitmap = 51'b111111111111110000000000000000000000000000000000000;
        12'b010010011001: bitmap = 51'b111111111111111000000000000000000000000000000000000;
        12'b010010011010: bitmap = 51'b111111111111111000000000000000000000000000000000000;
        12'b010010011011: bitmap = 51'b111111111111111100000000000000000000000000000000000;
        12'b010010011100: bitmap = 51'b111111111111111100000000000000000000000000000000000;
        12'b010010011101: bitmap = 51'b111111111111111110000000000000000000000000000000000;
        12'b010010011110: bitmap = 51'b111111111111111110000000000000000000000000000000000;
        12'b010010011111: bitmap = 51'b111111111111111111000000000000000000000000000000000;
        12'b010010100000: bitmap = 51'b111111111111111111100000000000000000000000000000000;
        12'b010010100001: bitmap = 51'b111111111111111111110000000000000000000000000000000;
        12'b010010100010: bitmap = 51'b111111111111111111111000000000000000000000000000000;
        12'b010010100011: bitmap = 51'b111111111111111111111110000000000000000000000000000;
        12'b010010100100: bitmap = 51'b111111111111111111111111100000000000000000000000000;
        12'b010010100101: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b010010100110: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b010010100111: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b010010101000: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b010010101001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b010010101010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b010010101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b010010101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b010010101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b010010101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b010010101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b010010110000: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b010010110001: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b010010110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b010010110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b010010110100: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b010010110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b010010110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b010010110111: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b010010111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b010010111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b010010111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b010010111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;

        
        12'b010011000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b010011000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b010011000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b010011000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b010011000100: bitmap = 51'b000000000000000000011111111111110000000000000000000;
        12'b010011000101: bitmap = 51'b000000000000000011111111111111100000000000000000000;
        12'b010011000110: bitmap = 51'b000000000000001111111111111111100000000000000000000;
        12'b010011000111: bitmap = 51'b000000000000011111111111111111000000000000000000000;
        12'b010011001000: bitmap = 51'b000000000001111111111111111111000000000000000000000;
        12'b010011001001: bitmap = 51'b000000000111111111111111111110000000000000000000000;
        12'b010011001010: bitmap = 51'b000000001111111111111111111110000000000000000000000;
        12'b010011001011: bitmap = 51'b000000111111111111111111111100000000000000011000000;
        12'b010011001100: bitmap = 51'b000011111111111111111111111000000000000000011110000;
        12'b010011001101: bitmap = 51'b000111111111111111111111111000000000000000111111000;
        12'b010011001110: bitmap = 51'b011111111111111111111111110000000000000000111111110;
        12'b010011001111: bitmap = 51'b111111111111111111111111110000000000000001111111111;
        12'b010011010000: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b010011010001: bitmap = 51'b111111111111111111111111100000000000000011111111111;
        12'b010011010010: bitmap = 51'b111111111111111111111111000000000000000011111111111;
        12'b010011010011: bitmap = 51'b111111111111111111111110000000000000000111111111111;
        12'b010011010100: bitmap = 51'b111111111111111111111110000000000000001111111111111;
        12'b010011010101: bitmap = 51'b111111111111111111111100000000000000001111111111111;
        12'b010011010110: bitmap = 51'b111111111111111111111100000000000000011111111111111;
        12'b010011010111: bitmap = 51'b111111111111111111111000000000000000000000000000000;
        12'b010011011000: bitmap = 51'b111111111111111111111000000000000000000000000000000;
        12'b010011011001: bitmap = 51'b111111111111111111110000000000000000000000000000000;
        12'b010011011010: bitmap = 51'b111111111111111111110000000000000000000000000000000;
        12'b010011011011: bitmap = 51'b111111111111111111100000000000000000000000000000000;
        12'b010011011100: bitmap = 51'b111111111111111111100000000000000000000000000000000;
        12'b010011011101: bitmap = 51'b111111111111111111100000000000000000000000000000000;
        12'b010011011110: bitmap = 51'b111111111111111111100000000000000000000000000000000;
        12'b010011011111: bitmap = 51'b111111111111111111100000000000000000000000000000000;
        12'b010011100000: bitmap = 51'b111111111111111111100000000000000000000000000000000;
        12'b010011100001: bitmap = 51'b111111111111111111110000000000000000000000000000000;
        12'b010011100010: bitmap = 51'b111111111111111111110000000000000000000000000000000;
        12'b010011100011: bitmap = 51'b111111111111111111111000000000000000000000000000000;
        12'b010011100100: bitmap = 51'b111111111111111111111000000000000000000000000000000;
        12'b010011100101: bitmap = 51'b111111111111111111111100000000000000001111111111111;
        12'b010011100110: bitmap = 51'b111111111111111111111110000000000000001111111111111;
        12'b010011100111: bitmap = 51'b111111111111111111111110000000000000000111111111111;
        12'b010011101000: bitmap = 51'b111111111111111111111111000000000000000111111111111;
        12'b010011101001: bitmap = 51'b111111111111111111111111000000000000000011111111111;
        12'b010011101010: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b010011101011: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b010011101100: bitmap = 51'b111111111111111111111111110000000000000000111111111;
        12'b010011101101: bitmap = 51'b011111111111111111111111110000000000000000111111110;
        12'b010011101110: bitmap = 51'b000111111111111111111111111000000000000000011111000;
        12'b010011101111: bitmap = 51'b000011111111111111111111111100000000000000011110000;
        12'b010011110000: bitmap = 51'b000000111111111111111111111100000000000000001000000;
        12'b010011110001: bitmap = 51'b000000001111111111111111111110000000000000000000000;
        12'b010011110010: bitmap = 51'b000000000111111111111111111110000000000000000000000;
        12'b010011110011: bitmap = 51'b000000000001111111111111111111000000000000000000000;
        12'b010011110100: bitmap = 51'b000000000000011111111111111111000000000000000000000;
        12'b010011110101: bitmap = 51'b000000000000001111111111111111100000000000000000000;
        12'b010011110110: bitmap = 51'b000000000000000011111111111111100000000000000000000;
        12'b010011110111: bitmap = 51'b000000000000000000011111111111110000000000000000000;
        12'b010011111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b010011111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b010011111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b010011111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        
        //shape 3
        12'b011000000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b011000000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b011000000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b011000000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b011000000100: bitmap = 51'b000000000000000000011111111111111000000000000000000;
        12'b011000000101: bitmap = 51'b000000000000000000001111111111111110000000000000000;
        12'b011000000110: bitmap = 51'b000000000000000000001111111111111111100000000000000;
        12'b011000000111: bitmap = 51'b000000000000000000000111111111111111110000000000000;
        12'b011000001000: bitmap = 51'b000000000000000000000011111111111111111100000000000;
        12'b011000001001: bitmap = 51'b000000000000000000000001111111111111111111000000000;
        12'b011000001010: bitmap = 51'b000000000000000000000001111111111111111111100000000;
        12'b011000001011: bitmap = 51'b000000100000000000000000111111111111111111111000000;
        12'b011000001100: bitmap = 51'b000011110000000000000000011111111111111111111110000;
        12'b011000001101: bitmap = 51'b000111111000000000000000011111111111111111111111000;
        12'b011000001110: bitmap = 51'b011111111000000000000000011111111111111111111111110;
        12'b011000001111: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b011000010000: bitmap = 51'b111111111110000000000000001111111111111111111111111;
        12'b011000010001: bitmap = 51'b111111111111000000000000000111111111111111111111111;
        12'b011000010010: bitmap = 51'b111111111111000000000000000111111111111111111111111;
        12'b011000010011: bitmap = 51'b111111111111000000000000000011111111111111111111111;
        12'b011000010100: bitmap = 51'b111111111111100000000000000011111111111111111111111;
        12'b011000010101: bitmap = 51'b111111111111110000000000000001111111111111111111111;
        12'b011000010110: bitmap = 51'b111111111111110000000000000001111111111111111111111;
        12'b011000010111: bitmap = 51'b111111111111100000000000000001111111111111111111111;
        12'b011000011000: bitmap = 51'b111111111111000000000000000001111111111111111111111;
        12'b011000011001: bitmap = 51'b000000000000000000000000000000111111111111111111111;
        12'b011000011010: bitmap = 51'b000000000000000000000000000000111111111111111111111;
        12'b011000011011: bitmap = 51'b000000000000000000000000000000111111111111111111111;
        12'b011000011100: bitmap = 51'b000000000000000000000000000000111111111111111111111;
        12'b011000011101: bitmap = 51'b000000000000000000000000000000111111111111111111111;
        12'b011000011110: bitmap = 51'b000000000000000000000000000001111111111111111111111;
        12'b011000011111: bitmap = 51'b000000000000000000000000000011111111111111111111111;
        12'b011000100000: bitmap = 51'b000000000000000000000000000111111111111111111111111;
        12'b011000100001: bitmap = 51'b000000000000000000000000111111111111111111111111111;
        12'b011000100010: bitmap = 51'b000000000000000000000111111111111111111111111111111;
        12'b011000100011: bitmap = 51'b000000000000000000111111111111111111111111111111111;
        12'b011000100100: bitmap = 51'b000000000000011111111111111111111111111111111111111;
        12'b011000100101: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011000100110: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011000100111: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011000101000: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011000101001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011000101010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011000101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011000101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011000101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b011000101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b011000101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b011000110000: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b011000110001: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b011000110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b011000110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b011000110100: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b011000110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b011000110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b011000110111: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b011000111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b011000111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b011000111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b011000111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        
        12'b011001000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b011001000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b011001000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b011001000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b011001000100: bitmap = 51'b000000000000000000011111111111110000000000000000000;
        12'b011001000101: bitmap = 51'b000000000000000000001111111111110000000000000000000;
        12'b011001000110: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b011001000111: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b011001001000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b011001001001: bitmap = 51'b000000000000000000000111111111100000000000000000000;
        12'b011001001010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b011001001011: bitmap = 51'b000000100000000000000111111111000000000000001000000;
        12'b011001001100: bitmap = 51'b000011100000000000000011111111000000000000011110000;
        12'b011001001101: bitmap = 51'b000111110000000000000001111110000000000000011111000;
        12'b011001001110: bitmap = 51'b011111110000000000000000111100000000000000111111110;
        12'b011001001111: bitmap = 51'b111111111000000000000000011000000000000000111111111;
        12'b011001010000: bitmap = 51'b111111111000000000000000000000000000000000111111111;
        12'b011001010001: bitmap = 51'b111111111100000000000000000000000000000001111111111;
        12'b011001010010: bitmap = 51'b111111111100000000000000000000000000000001111111111;
        12'b011001010011: bitmap = 51'b111111111100000000000000000000000000000011111111111;
        12'b011001010100: bitmap = 51'b111111111110000000000000000000000000000011111111111;
        12'b011001010101: bitmap = 51'b111111111110000000000000000000000000000011111111111;
        12'b011001010110: bitmap = 51'b111111111111000000000000000000000000000111111111111;
        12'b011001010111: bitmap = 51'b111111111111100000000000000000000000001111111111111;
        12'b011001011000: bitmap = 51'b111111111111110000000000000000000000001111111111111;
        12'b011001011001: bitmap = 51'b111111111111110000000000000000000000011111111111111;
        12'b011001011010: bitmap = 51'b111111111111111000000000000000000000111111111111111;
        12'b011001011011: bitmap = 51'b111111111111111100000000000000000001111111111111111;
        12'b011001011100: bitmap = 51'b111111111111111110000000000000000011111111111111111;
        12'b011001011101: bitmap = 51'b111111111111111111000000000000000111111111111111111;
        12'b011001011110: bitmap = 51'b111111111111111111100000000000001111111111111111111;
        12'b011001011111: bitmap = 51'b111111111111111111110000000000011111111111111111111;
        12'b011001100000: bitmap = 51'b111111111111111111111000000000111111111111111111111;
        12'b011001100001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011001100010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011001100011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011001100100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011001100101: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011001100110: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011001100111: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011001101000: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011001101001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011001101010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011001101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011001101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011001101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b011001101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b011001101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b011001110000: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b011001110001: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b011001110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b011001110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b011001110100: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b011001110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b011001110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b011001110111: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b011001111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b011001111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b011001111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b011001111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        
        12'b011010000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b011010000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b011010000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b011010000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b011010000100: bitmap = 51'b000000000000000000111111111111110000000000000000000;
        12'b011010000101: bitmap = 51'b000000000000000011111111111111100000000000000000000;
        12'b011010000110: bitmap = 51'b000000000000001111111111111111100000000000000000000;
        12'b011010000111: bitmap = 51'b000000000000011111111111111111000000000000000000000;
        12'b011010001000: bitmap = 51'b000000000001111111111111111110000000000000000000000;
        12'b011010001001: bitmap = 51'b000000000111111111111111111100000000000000000000000;
        12'b011010001010: bitmap = 51'b000000001111111111111111111100000000000000000000000;
        12'b011010001011: bitmap = 51'b000000111111111111111111111000000000000000001000000;
        12'b011010001100: bitmap = 51'b000011111111111111111111110000000000000000011110000;
        12'b011010001101: bitmap = 51'b000111111111111111111111110000000000000000111111000;
        12'b011010001110: bitmap = 51'b011111111111111111111111110000000000000000111111110;
        12'b011010001111: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b011010010000: bitmap = 51'b111111111111111111111111100000000000000011111111111;
        12'b011010010001: bitmap = 51'b111111111111111111111111000000000000000111111111111;
        12'b011010010010: bitmap = 51'b111111111111111111111111000000000000000111111111111;
        12'b011010010011: bitmap = 51'b111111111111111111111110000000000000000111111111111;
        12'b011010010100: bitmap = 51'b111111111111111111111110000000000000001111111111111;
        12'b011010010101: bitmap = 51'b111111111111111111111100000000000000011111111111111;
        12'b011010010110: bitmap = 51'b111111111111111111111100000000000000011111111111111;
        12'b011010010111: bitmap = 51'b111111111111111111111100000000000000001111111111111;
        12'b011010011000: bitmap = 51'b111111111111111111111100000000000000000111111111111;
        12'b011010011001: bitmap = 51'b111111111111111111111000000000000000000000000000000;
        12'b011010011010: bitmap = 51'b111111111111111111111000000000000000000000000000000;
        12'b011010011011: bitmap = 51'b111111111111111111111000000000000000000000000000000;
        12'b011010011100: bitmap = 51'b111111111111111111111000000000000000000000000000000;
        12'b011010011101: bitmap = 51'b111111111111111111111000000000000000000000000000000;
        12'b011010011110: bitmap = 51'b111111111111111111111100000000000000000000000000000;
        12'b011010011111: bitmap = 51'b111111111111111111111110000000000000000000000000000;
        12'b011010100000: bitmap = 51'b111111111111111111111111000000000000000000000000000;
        12'b011010100001: bitmap = 51'b111111111111111111111111111000000000000000000000000;
        12'b011010100010: bitmap = 51'b111111111111111111111111111111000000000000000000000;
        12'b011010100011: bitmap = 51'b111111111111111111111111111111111000000000000000000;
        12'b011010100100: bitmap = 51'b111111111111111111111111111111111111110000000000000;
        12'b011010100101: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011010100110: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011010100111: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011010101000: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011010101001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011010101010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011010101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011010101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b011010101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b011010101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b011010101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b011010110000: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b011010110001: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b011010110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b011010110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b011010110100: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b011010110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b011010110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b011010110111: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b011010111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b011010111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b011010111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b011010111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;

       //shape 4
        12'b100000000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b100000000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b100000000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b100000000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b100000000100: bitmap = 51'b000000000000000000011111111111110000000000000000000;
        12'b100000000101: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b100000000110: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b100000000111: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b100000001000: bitmap = 51'b000000000000000000000011111111000000000000000000000;
        12'b100000001001: bitmap = 51'b000000000000000000000001111110000000000000000000000;
        12'b100000001010: bitmap = 51'b000000000000000000000001111110000000000000000000000;
        12'b100000001011: bitmap = 51'b000000100000000000000000111100000000000000001000000;
        12'b100000001100: bitmap = 51'b000011110000000000000000011000000000000000011110000;
        12'b100000001101: bitmap = 51'b000111111000000000000000001000000000000000011111000;
        12'b100000001110: bitmap = 51'b011111111000000000000000000000000000000000111111110;
        12'b100000001111: bitmap = 51'b111111111100000000000000000000000000000000111111111;
        12'b100000010000: bitmap = 51'b111111111110000000000000000000000000000001111111111;
        12'b100000010001: bitmap = 51'b111111111111000000000000000000000000000001111111111;
        12'b100000010010: bitmap = 51'b111111111111000000000000000000000000000011111111111;
        12'b100000010011: bitmap = 51'b111111111111000000000000000000000000000111111111111;
        12'b100000010100: bitmap = 51'b111111111111100000000000000000000000000111111111111;
        12'b100000010101: bitmap = 51'b111111111111100000000000000000000000001111111111111;
        12'b100000010110: bitmap = 51'b111111111111100000000000000000000000001111111111111;
        12'b100000010111: bitmap = 51'b111111111111100000000000000000000000011111111111111;
        12'b100000011000: bitmap = 51'b111111111111000000000000000000000000011111111111111;
        12'b100000011001: bitmap = 51'b000000000000000000000000000000000000111111111111111;
        12'b100000011010: bitmap = 51'b000000000000000000000000000000000001111111111111111;
        12'b100000011011: bitmap = 51'b000000000000000000000000000000000001111111111111111;
        12'b100000011100: bitmap = 51'b000000000000000000000000000000000011111111111111111;
        12'b100000011101: bitmap = 51'b000000000000000000000000000000000011111111111111111;
        12'b100000011110: bitmap = 51'b000000000000000000000000000000000111111111111111111;
        12'b100000011111: bitmap = 51'b000000000000000000000000000000000111111111111111111;
        12'b100000100000: bitmap = 51'b000000000000000000000000000000001111111111111111111;
        12'b100000100001: bitmap = 51'b000000000000000000000000000000001111111111111111111;
        12'b100000100010: bitmap = 51'b000000000000000000000000000000011111111111111111111;
        12'b100000100011: bitmap = 51'b000000000000000000000000000000111111111111111111111;
        12'b100000100100: bitmap = 51'b000000000000000000000000000000111111111111111111111;
        12'b100000100101: bitmap = 51'b111111111111100000000000000001111111111111111111111;
        12'b100000100110: bitmap = 51'b111111111111100000000000000001111111111111111111111;
        12'b100000100111: bitmap = 51'b111111111111000000000000000011111111111111111111111;
        12'b100000101000: bitmap = 51'b111111111111000000000000000011111111111111111111111;
        12'b100000101001: bitmap = 51'b111111111110000000000000000111111111111111111111111;
        12'b100000101010: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b100000101011: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b100000101100: bitmap = 51'b111111111000000000000000011111111111111111111111111;
        12'b100000101101: bitmap = 51'b011111111000000000000000011111111111111111111111110;
        12'b100000101110: bitmap = 51'b000111110000000000000000111111111111111111111111000;
        12'b100000101111: bitmap = 51'b000011110000000000000000111111111111111111111110000;
        12'b100000110000: bitmap = 51'b000000100000000000000001111111111111111111111000000;
        12'b100000110001: bitmap = 51'b000000000000000000000011111111111111111111100000000;
        12'b100000110010: bitmap = 51'b000000000000000000000011111111111111111111000000000;
        12'b100000110011: bitmap = 51'b000000000000000000000111111111111111111100000000000;
        12'b100000110100: bitmap = 51'b000000000000000000000111111111111111110000000000000;
        12'b100000110101: bitmap = 51'b000000000000000000001111111111111111100000000000000;
        12'b100000110110: bitmap = 51'b000000000000000000001111111111111110000000000000000;
        12'b100000110111: bitmap = 51'b000000000000000000011111111111111000000000000000000;
        12'b100000111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b100000111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b100000111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b100000111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;

        12'b100001000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b100001000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b100001000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b100001000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b100001000100: bitmap = 51'b000000000000000000011111111111110000000000000000000;
        12'b100001000101: bitmap = 51'b000000000000000000001111111111110000000000000000000;
        12'b100001000110: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b100001000111: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b100001001000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b100001001001: bitmap = 51'b000000000000000000000111111111100000000000000000000;
        12'b100001001010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b100001001011: bitmap = 51'b000000100000000000000111111111000000000000001000000;
        12'b100001001100: bitmap = 51'b000011100000000000000011111111000000000000011110000;
        12'b100001001101: bitmap = 51'b000111110000000000000001111110000000000000011111000;
        12'b100001001110: bitmap = 51'b011111110000000000000000111100000000000000111111110;
        12'b100001001111: bitmap = 51'b111111111000000000000000011000000000000000111111111;
        12'b100001010000: bitmap = 51'b111111111000000000000000000000000000000000111111111;
        12'b100001010001: bitmap = 51'b111111111100000000000000000000000000000001111111111;
        12'b100001010010: bitmap = 51'b111111111100000000000000000000000000000001111111111;
        12'b100001010011: bitmap = 51'b111111111100000000000000000000000000000011111111111;
        12'b100001010100: bitmap = 51'b111111111110000000000000000000000000000011111111111;
        12'b100001010101: bitmap = 51'b111111111110000000000000000000000000000011111111111;
        12'b100001010110: bitmap = 51'b111111111111000000000000000000000000000111111111111;
        12'b100001010111: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b100001011000: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b100001011001: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b100001011010: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b100001011011: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b100001011100: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b100001011101: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b100001011110: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b100001011111: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b100001100000: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b100001100001: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b100001100010: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b100001100011: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b100001100100: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b100001100101: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b100001100110: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b100001100111: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b100001101000: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b100001101001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b100001101010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b100001101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b100001101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b100001101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b100001101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b100001101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b100001110000: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b100001110001: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b100001110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b100001110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b100001110100: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b100001110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b100001110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b100001110111: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b100001111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b100001111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b100001111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b100001111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;

        12'b100010000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b100010000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b100010000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b100010000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b100010000100: bitmap = 51'b000000000000000000011111111111110000000000000000000;
        12'b100010000101: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b100010000110: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b100010000111: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b100010001000: bitmap = 51'b000000000000000000000111111110000000000000000000000;
        12'b100010001001: bitmap = 51'b000000000000000000000011111100000000000000000000000;
        12'b100010001010: bitmap = 51'b000000000000000000000011111100000000000000000000000;
        12'b100010001011: bitmap = 51'b000000100000000000000001111000000000000000001000000;
        12'b100010001100: bitmap = 51'b000011110000000000000000110000000000000000011110000;
        12'b100010001101: bitmap = 51'b000111110000000000000000100000000000000000111111000;
        12'b100010001110: bitmap = 51'b011111111000000000000000000000000000000000111111110;
        12'b100010001111: bitmap = 51'b111111111000000000000000000000000000000001111111111;
        12'b100010010000: bitmap = 51'b111111111100000000000000000000000000000011111111111;
        12'b100010010001: bitmap = 51'b111111111100000000000000000000000000000111111111111;
        12'b100010010010: bitmap = 51'b111111111110000000000000000000000000000111111111111;
        12'b100010010011: bitmap = 51'b111111111111000000000000000000000000000111111111111;
        12'b100010010100: bitmap = 51'b111111111111000000000000000000000000001111111111111;
        12'b100010010101: bitmap = 51'b111111111111100000000000000000000000001111111111111;
        12'b100010010110: bitmap = 51'b111111111111100000000000000000000000001111111111111;
        12'b100010010111: bitmap = 51'b111111111111110000000000000000000000001111111111111;
        12'b100010011000: bitmap = 51'b111111111111110000000000000000000000000111111111111;
        12'b100010011001: bitmap = 51'b111111111111111000000000000000000000000000000000000;
        12'b100010011010: bitmap = 51'b111111111111111100000000000000000000000000000000000;
        12'b100010011011: bitmap = 51'b111111111111111100000000000000000000000000000000000;
        12'b100010011100: bitmap = 51'b111111111111111110000000000000000000000000000000000;
        12'b100010011101: bitmap = 51'b111111111111111110000000000000000000000000000000000;
        12'b100010011110: bitmap = 51'b111111111111111111000000000000000000000000000000000;
        12'b100010011111: bitmap = 51'b111111111111111111000000000000000000000000000000000;
        12'b100010100000: bitmap = 51'b111111111111111111100000000000000000000000000000000;
        12'b100010100001: bitmap = 51'b111111111111111111100000000000000000000000000000000;
        12'b100010100010: bitmap = 51'b111111111111111111110000000000000000000000000000000;
        12'b100010100011: bitmap = 51'b111111111111111111111000000000000000000000000000000;
        12'b100010100100: bitmap = 51'b111111111111111111111000000000000000000000000000000;
        12'b100010100101: bitmap = 51'b111111111111111111111100000000000000001111111111111;
        12'b100010100110: bitmap = 51'b111111111111111111111100000000000000001111111111111;
        12'b100010100111: bitmap = 51'b111111111111111111111110000000000000000111111111111;
        12'b100010101000: bitmap = 51'b111111111111111111111110000000000000000111111111111;
        12'b100010101001: bitmap = 51'b111111111111111111111111000000000000000011111111111;
        12'b100010101010: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b100010101011: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b100010101100: bitmap = 51'b111111111111111111111111110000000000000000111111111;
        12'b100010101101: bitmap = 51'b011111111111111111111111110000000000000000111111110;
        12'b100010101110: bitmap = 51'b000111111111111111111111111000000000000000011111000;
        12'b100010101111: bitmap = 51'b000011111111111111111111111000000000000000011110000;
        12'b100010110000: bitmap = 51'b000000111111111111111111111100000000000000001000000;
        12'b100010110001: bitmap = 51'b000000001111111111111111111110000000000000000000000;
        12'b100010110010: bitmap = 51'b000000000111111111111111111110000000000000000000000;
        12'b100010110011: bitmap = 51'b000000000001111111111111111111000000000000000000000;
        12'b100010110100: bitmap = 51'b000000000000011111111111111111000000000000000000000;
        12'b100010110101: bitmap = 51'b000000000000001111111111111111100000000000000000000;
        12'b100010110110: bitmap = 51'b000000000000000011111111111111100000000000000000000;
        12'b100010110111: bitmap = 51'b000000000000000000111111111111110000000000000000000;
        12'b100010111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b100010111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b100010111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b100010111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        
      //shape 5
         12'b101000000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b101000000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b101000000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b101000000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b101000000100: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b101000000101: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b101000000110: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b101000000111: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b101000001000: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b101000001001: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b101000001010: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b101000001011: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b101000001100: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b101000001101: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b101000001110: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b101000001111: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101000010000: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101000010001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101000010010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101000010011: bitmap = 51'b111111111111111111111100000001111111111111111111111;
        12'b101000010100: bitmap = 51'b111111111111111111110000000000011111111111111111111;
        12'b101000010101: bitmap = 51'b111111111111111111100000000000001111111111111111111;
        12'b101000010110: bitmap = 51'b111111111111111110000000000000000011111111111111111;
        12'b101000010111: bitmap = 51'b000000000000000000000000000000000011111111111111111;
        12'b101000011000: bitmap = 51'b000000000000000000000000000000000000101111111111111;
        12'b101000011001: bitmap = 51'b000000000000000000000000000000000000111111111111111;
        12'b101000011010: bitmap = 51'b000000000000000000000000000000000000111111111111111;
        12'b101000011011: bitmap = 51'b000000000000000000000000000000000000011111111111111;
        12'b101000011100: bitmap = 51'b000000000000000000000000000000000000011111111111111;
        12'b101000011101: bitmap = 51'b000000000000000000000000000000000000011111111111111;
        12'b101000011110: bitmap = 51'b000000000000000000000000000000000000011111111111111;
        12'b101000011111: bitmap = 51'b000000000000000000000000000000000000011111111111111;
        12'b101000100000: bitmap = 51'b000000000000000000000000000000000000011111111111111;
        12'b101000100001: bitmap = 51'b000000000000000000000000000000000000111111111111111;
        12'b101000100010: bitmap = 51'b000000000000000000000000000000000000111111111111111;
        12'b101000100011: bitmap = 51'b000000000000000000000000000000000001111111111111111;
        12'b101000100100: bitmap = 51'b000000000000000000000000000000000011111111111111111;
        12'b101000100101: bitmap = 51'b111111111111111110000000000000000011111111111111111;
        12'b101000100110: bitmap = 51'b111111111111111111100000000000001111111111111111111;
        12'b101000100111: bitmap = 51'b111111111111111111110000000000011111111111111111111;
        12'b101000101000: bitmap = 51'b111111111111111111111100000001111111111111111111111;
        12'b101000101001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101000101010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101000101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101000101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101000101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b101000101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b101000101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b101000110000: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b101000110001: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b101000110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b101000110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b101000110100: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b101000110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b101000110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b101000110111: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b101000111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b101000111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b101000111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b101000111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        
        
        
        12'b101001000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b101001000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b101001000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b101001000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b101001000100: bitmap = 51'b000000000000000000011111111111111000000000000000000;
        12'b101001000101: bitmap = 51'b000000000000000000001111111111111110000000000000000;
        12'b101001000110: bitmap = 51'b000000000000000000001111111111111111100000000000000;
        12'b101001000111: bitmap = 51'b000000000000000000000111111111111111110000000000000;
        12'b101001001000: bitmap = 51'b000000000000000000000111111111111111111100000000000;
        12'b101001001001: bitmap = 51'b000000000000000000000011111111111111111111000000000;
        12'b101001001010: bitmap = 51'b000000000000000000000011111111111111111111100000000;
        12'b101001001011: bitmap = 51'b000000100000000000000001111111111111111111111000000;
        12'b101001001100: bitmap = 51'b000011110000000000000000111111111111111111111110000;
        12'b101001001101: bitmap = 51'b000111110000000000000000111111111111111111111111000;
        12'b101001001110: bitmap = 51'b011111111000000000000000011111111111111111111111110;
        12'b101001001111: bitmap = 51'b111111111000000000000000011111111111111111111111111;
        12'b101001010000: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b101001010001: bitmap = 51'b111111111100000000000000000111111111111111111111111;
        12'b101001010010: bitmap = 51'b111111111110000000000000000011111111111111111111111;
        12'b101001010011: bitmap = 51'b111111111110000000000000000000001111111111111111111;
        12'b101001010100: bitmap = 51'b111111111111000000000000000000000011111111111111111;
        12'b101001010101: bitmap = 51'b111111111111100000000000000000000001111111111111111;
        12'b101001010110: bitmap = 51'b111111111111100000000000000000000000111111111111111;
        12'b101001010111: bitmap = 51'b111111111111110000000000000000000000011111111111111;
        12'b101001011000: bitmap = 51'b111111111111110000000000000000000000011111111111111;
        12'b101001011001: bitmap = 51'b111111111111111000000000000000000000001111111111111;
        12'b101001011010: bitmap = 51'b111111111111111000000000000000000000001111111111111;
        12'b101001011011: bitmap = 51'b111111111111111000000000000000000000000111111111111;
        12'b101001011100: bitmap = 51'b111111111111110000000000000000000000000111111111111;
        12'b101001011101: bitmap = 51'b111111111111110000000000000000000000000111111111111;
        12'b101001011110: bitmap = 51'b111111111111110000000000000000000000000111111111111;
        12'b101001011111: bitmap = 51'b111111111111110000000000000000000000000111111111111;
        12'b101001100000: bitmap = 51'b111111111111110000000000000000000000000111111111111;
        12'b101001100001: bitmap = 51'b111111111111110000000000000000000000000111111111111;
        12'b101001100010: bitmap = 51'b111111111111111000000000000000000000001111111111111;
        12'b101001100011: bitmap = 51'b111111111111111000000000000000000000001111111111111;
        12'b101001100100: bitmap = 51'b111111111111111100000000000000000000001111111111111;
        12'b101001100101: bitmap = 51'b111111111111111100000000000000000000011111111111111;
        12'b101001100110: bitmap = 51'b111111111111111110000000000000000000111111111111111;
        12'b101001100111: bitmap = 51'b111111111111111111000000000000000001111111111111111;
        12'b101001101000: bitmap = 51'b111111111111111111100000000000000011111111111111111;
        12'b101001101001: bitmap = 51'b111111111111111111111000000000001111111111111111111;
        12'b101001101010: bitmap = 51'b111111111111111111111110000000111111111111111111111;
        12'b101001101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101001101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101001101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b101001101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b101001101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b101001110000: bitmap = 51'b000000111111111111111111111111111111111111111100000;
        12'b101001110001: bitmap = 51'b000000001111111111111111111111111111111111110000000;
        12'b101001110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b101001110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b101001110100: bitmap = 51'b000000000000011111111111111111111111111000000000000;
        12'b101001110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b101001110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b101001110111: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b101001111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b101001111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b101001111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b101001111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        
        12'b101010000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b101010000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b101010000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b101010000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b101010000100: bitmap = 51'b000000000000000000111111111111110000000000000000000;
        12'b101010000101: bitmap = 51'b000000000000000011111111111111100000000000000000000;
        12'b101010000110: bitmap = 51'b000000000000001111111111111111100000000000000000000;
        12'b101010000111: bitmap = 51'b000000000000011111111111111111000000000000000000000;
        12'b101010001000: bitmap = 51'b000000000001111111111111111111000000000000000000000;
        12'b101010001001: bitmap = 51'b000000000111111111111111111110000000000000000000000;
        12'b101010001010: bitmap = 51'b000000001111111111111111111110000000000000000000000;
        12'b101010001011: bitmap = 51'b000000111111111111111111111100000000000000001000000;
        12'b101010001100: bitmap = 51'b000011111111111111111111111000000000000000011110000;
        12'b101010001101: bitmap = 51'b000111111111111111111111111000000000000000011111000;
        12'b101010001110: bitmap = 51'b011111111111111111111111110000000000000000111111110;
        12'b101010001111: bitmap = 51'b111111111111111111111111110000000000000000111111111;
        12'b101010010000: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b101010010001: bitmap = 51'b111111111111111111111111000000000000000001111111111;
        12'b101010010010: bitmap = 51'b111111111111111111111110000000000000000011111111111;
        12'b101010010011: bitmap = 51'b111111111111111111100000000000000000000011111111111;
        12'b101010010100: bitmap = 51'b111111111111111110000000000000000000000111111111111;
        12'b101010010101: bitmap = 51'b111111111111111100000000000000000000001111111111111;
        12'b101010010110: bitmap = 51'b111111111111111000000000000000000000001111111111111;
        12'b101010010111: bitmap = 51'b111111111111110000000000000000000000011111111111111;
        12'b101010011000: bitmap = 51'b111111111111110000000000000000000000011111111111111;
        12'b101010011001: bitmap = 51'b111111111111100000000000000000000000111111111111111;
        12'b101010011010: bitmap = 51'b111111111111100000000000000000000000111111111111111;
        12'b101010011011: bitmap = 51'b111111111111000000000000000000000000111111111111111;
        12'b101010011100: bitmap = 51'b111111111111000000000000000000000000011111111111111;
        12'b101010011101: bitmap = 51'b111111111111000000000000000000000000011111111111111;
        12'b101010011110: bitmap = 51'b111111111111000000000000000000000000011111111111111;
        12'b101010011111: bitmap = 51'b111111111111000000000000000000000000011111111111111;
        12'b101010100000: bitmap = 51'b111111111111000000000000000000000000011111111111111;
        12'b101010100001: bitmap = 51'b111111111111000000000000000000000000011111111111111;
        12'b101010100010: bitmap = 51'b111111111111100000000000000000000000111111111111111;
        12'b101010100011: bitmap = 51'b111111111111100000000000000000000000111111111111111;
        12'b101010100100: bitmap = 51'b111111111111100000000000000000000001111111111111111;
        12'b101010100101: bitmap = 51'b111111111111110000000000000000000001111111111111111;
        12'b101010100110: bitmap = 51'b111111111111111000000000000000000011111111111111111;
        12'b101010100111: bitmap = 51'b111111111111111100000000000000000111111111111111111;
        12'b101010101000: bitmap = 51'b111111111111111110000000000000001111111111111111111;
        12'b101010101001: bitmap = 51'b111111111111111111100000000000111111111111111111111;
        12'b101010101010: bitmap = 51'b111111111111111111111000000011111111111111111111111;
        12'b101010101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101010101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101010101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b101010101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b101010101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b101010110000: bitmap = 51'b000001111111111111111111111111111111111111111000000;
        12'b101010110001: bitmap = 51'b000000011111111111111111111111111111111111100000000;
        12'b101010110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b101010110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b101010110100: bitmap = 51'b000000000000111111111111111111111111110000000000000;
        12'b101010110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b101010110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b101010110111: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b101010111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b101010111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b101010111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b101010111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        
        12'b101011000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b101011000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b101011000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b101011000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b101011000100: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b101011000101: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b101011000110: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b101011000111: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b101011001000: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b101011001001: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b101011001010: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b101011001011: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b101011001100: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b101011001101: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b101011001110: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b101011001111: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101011010000: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101011010001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101011010010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101011010011: bitmap = 51'b111111111111111111111100000001111111111111111111111;
        12'b101011010100: bitmap = 51'b111111111111111111110000000000011111111111111111111;
        12'b101011010101: bitmap = 51'b111111111111111111100000000000001111111111111111111;
        12'b101011010110: bitmap = 51'b111111111111111110000000000000000011111111111111111;
        12'b101011010111: bitmap = 51'b111111111111111110000000000000000000000000000000000;
        12'b101011011000: bitmap = 51'b111111111111101000000000000000000000000000000000000;
        12'b101011011001: bitmap = 51'b111111111111111000000000000000000000000000000000000;
        12'b101011011010: bitmap = 51'b111111111111111000000000000000000000000000000000000;
        12'b101011011011: bitmap = 51'b111111111111110000000000000000000000000000000000000;
        12'b101011011100: bitmap = 51'b111111111111110000000000000000000000000000000000000;
        12'b101011011101: bitmap = 51'b111111111111110000000000000000000000000000000000000;
        12'b101011011110: bitmap = 51'b111111111111110000000000000000000000000000000000000;
        12'b101011011111: bitmap = 51'b111111111111110000000000000000000000000000000000000;
        12'b101011100000: bitmap = 51'b111111111111110000000000000000000000000000000000000;
        12'b101011100001: bitmap = 51'b111111111111111000000000000000000000000000000000000;
        12'b101011100010: bitmap = 51'b111111111111111000000000000000000000000000000000000;
        12'b101011100011: bitmap = 51'b111111111111111100000000000000000000000000000000000;
        12'b101011100100: bitmap = 51'b111111111111111110000000000000000000000000000000000;
        12'b101011100101: bitmap = 51'b111111111111111110000000000000000011111111111111111;
        12'b101011100110: bitmap = 51'b111111111111111111100000000000001111111111111111111;
        12'b101011100111: bitmap = 51'b111111111111111111110000000000011111111111111111111;
        12'b101011101000: bitmap = 51'b111111111111111111111100000001111111111111111111111;
        12'b101011101001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101011101010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101011101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101011101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b101011101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b101011101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b101011101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b101011110000: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b101011110001: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b101011110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b101011110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b101011110100: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b101011110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b101011110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b101011110111: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b101011111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b101011111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b101011111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b101011111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        

      //shape 6
        12'b110000000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b110000000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b110000000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b110000000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b110000000100: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b110000000101: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b110000000110: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b110000000111: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b110000001000: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b110000001001: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b110000001010: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b110000001011: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b110000001100: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b110000001101: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b110000001110: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b110000001111: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110000010000: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110000010001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110000010010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110000010011: bitmap = 51'b111111111111111111111100000001111111111111111111111;
        12'b110000010100: bitmap = 51'b111111111111111111110000000000011111111111111111111;
        12'b110000010101: bitmap = 51'b111111111111111111100000000000001111111111111111111;
        12'b110000010110: bitmap = 51'b111111111111111110000000000000000011111111111111111;
        12'b110000010111: bitmap = 51'b000000000000000000000000000000000011111111111111111;
        12'b110000011000: bitmap = 51'b000000000000000000000000000000000000101111111111111;
        12'b110000011001: bitmap = 51'b000000000000000000000000111100000000111111111111111;
        12'b110000011010: bitmap = 51'b000000000000000000000001111110000000111111111111111;
        12'b110000011011: bitmap = 51'b000000000000000000000011111111000000011111111111111;
        12'b110000011100: bitmap = 51'b000000000000000000000111111111100000011111111111111;
        12'b110000011101: bitmap = 51'b000000000000000000000111111111100000011111111111111;
        12'b110000011110: bitmap = 51'b000000000000000000000111111111100000011111111111111;
        12'b110000011111: bitmap = 51'b000000000000000000000111111111100000011111111111111;
        12'b110000100000: bitmap = 51'b000000000000000000000011111111000000011111111111111;
        12'b110000100001: bitmap = 51'b000000000000000000000001111110000000111111111111111;
        12'b110000100010: bitmap = 51'b000000000000000000000000111100000000111111111111111;
        12'b110000100011: bitmap = 51'b000000000000000000000000000000000001111111111111111;
        12'b110000100100: bitmap = 51'b000000000000000000000000000000000011111111111111111;
        12'b110000100101: bitmap = 51'b111111111111111110000000000000000011111111111111111;
        12'b110000100110: bitmap = 51'b111111111111111111100000000000001111111111111111111;
        12'b110000100111: bitmap = 51'b111111111111111111110000000000011111111111111111111;
        12'b110000101000: bitmap = 51'b111111111111111111111100000001111111111111111111111;
        12'b110000101001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110000101010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110000101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110000101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110000101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b110000101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b110000101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b110000110000: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b110000110001: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b110000110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b110000110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b110000110100: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b110000110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b110000110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b110000110111: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b110000111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b110000111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b110000111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b110000111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        
        
        
        12'b110001000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b110001000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b110001000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b110001000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b110001000100: bitmap = 51'b000000000000000000011111111111111000000000000000000;
        12'b110001000101: bitmap = 51'b000000000000000000001111111111111110000000000000000;
        12'b110001000110: bitmap = 51'b000000000000000000000111111111111111100000000000000;
        12'b110001000111: bitmap = 51'b000000000000000000000111111111111111110000000000000;
        12'b110001001000: bitmap = 51'b000000000000000000000111111111111111111100000000000;
        12'b110001001001: bitmap = 51'b000000000000000000000011111111111111111111000000000;
        12'b110001001010: bitmap = 51'b000000000000000000000011111111111111111111100000000;
        12'b110001001011: bitmap = 51'b000000100000000000000001111111111111111111111000000;
        12'b110001001100: bitmap = 51'b000011100000000000000000111111111111111111111110000;
        12'b110001001101: bitmap = 51'b000111110000000000000000111111111111111111111111000;
        12'b110001001110: bitmap = 51'b011111111000000000000000011111111111111111111111110;
        12'b110001001111: bitmap = 51'b111111111100000000000000011111111111111111111111111;
        12'b110001010000: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b110001010001: bitmap = 51'b111111111110000000000000000111111111111111111111111;
        12'b110001010010: bitmap = 51'b111111111110000000000000000000111111111111111111111;
        12'b110001010011: bitmap = 51'b111111111111000000000000000000001111111111111111111;
        12'b110001010100: bitmap = 51'b111111111111000000000000000000000011111111111111111;
        12'b110001010101: bitmap = 51'b111111111111100000000000000000000001111111111111111;
        12'b110001010110: bitmap = 51'b111111111111100000000000000000000000111111111111111;
        12'b110001010111: bitmap = 51'b111111111111110000000000000000000000011111111111111;
        12'b110001011000: bitmap = 51'b111111111111110000000000000000000000011111111111111;
        12'b110001011001: bitmap = 51'b111111111111111000000000111110000000001111111111111;
        12'b110001011010: bitmap = 51'b111111111111111000000001111111000000001111111111111;
        12'b110001011011: bitmap = 51'b111111111111110000000011111111100000000111111111111;
        12'b110001011100: bitmap = 51'b111111111111110000000111111111110000000111111111111;
        12'b110001011101: bitmap = 51'b111111111111110000000111111111110000000111111111111;
        12'b110001011110: bitmap = 51'b111111111111110000000111111111110000000111111111111;
        12'b110001011111: bitmap = 51'b111111111111110000000111111111110000000111111111111;
        12'b110001100000: bitmap = 51'b111111111111110000000111111111110000000111111111111;
        12'b110001100001: bitmap = 51'b111111111111110000000011111111100000000111111111111;
        12'b110001100010: bitmap = 51'b111111111111111000000001111111000000001111111111111;
        12'b110001100011: bitmap = 51'b111111111111111000000000111110000000001111111111111;
        12'b110001100100: bitmap = 51'b111111111111111100000000000000000000001111111111111;
        12'b110001100101: bitmap = 51'b111111111111111100000000000000000000011111111111111;
        12'b110001100110: bitmap = 51'b111111111111111110000000000000000000111111111111111;
        12'b110001100111: bitmap = 51'b111111111111111111000000000000000001111111111111111;
        12'b110001101000: bitmap = 51'b111111111111111111100000000000000011111111111111111;
        12'b110001101001: bitmap = 51'b111111111111111111111000000000001111111111111111111;
        12'b110001101010: bitmap = 51'b111111111111111111111110000000111111111111111111111;
        12'b110001101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110001101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110001101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b110001101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b110001101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b110001110000: bitmap = 51'b000000111111111111111111111111111111111111111100000;
        12'b110001110001: bitmap = 51'b000000001111111111111111111111111111111111110000000;
        12'b110001110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b110001110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b110001110100: bitmap = 51'b000000000000011111111111111111111111111000000000000;
        12'b110001110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b110001110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b110001110111: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b110001111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b110001111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b110001111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b110001111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        
        12'b110010000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b110010000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b110010000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b110010000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b110010000100: bitmap = 51'b000000000000000000111111111111110000000000000000000;
        12'b110010000101: bitmap = 51'b000000000000000011111111111111100000000000000000000;
        12'b110010000110: bitmap = 51'b000000000000001111111111111111000000000000000000000;
        12'b110010000111: bitmap = 51'b000000000000011111111111111111000000000000000000000;
        12'b110010001000: bitmap = 51'b000000000001111111111111111111000000000000000000000;
        12'b110010001001: bitmap = 51'b000000000111111111111111111110000000000000000000000;
        12'b110010001010: bitmap = 51'b000000001111111111111111111110000000000000000000000;
        12'b110010001011: bitmap = 51'b000000111111111111111111111100000000000000001000000;
        12'b110010001100: bitmap = 51'b000011111111111111111111111000000000000000001110000;
        12'b110010001101: bitmap = 51'b000111111111111111111111111000000000000000011111000;
        12'b110010001110: bitmap = 51'b011111111111111111111111110000000000000000111111110;
        12'b110010001111: bitmap = 51'b111111111111111111111111110000000000000001111111111;
        12'b110010010000: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b110010010001: bitmap = 51'b111111111111111111111111000000000000000011111111111;
        12'b110010010010: bitmap = 51'b111111111111111111111000000000000000000011111111111;
        12'b110010010011: bitmap = 51'b111111111111111111100000000000000000000111111111111;
        12'b110010010100: bitmap = 51'b111111111111111110000000000000000000000111111111111;
        12'b110010010101: bitmap = 51'b111111111111111100000000000000000000001111111111111;
        12'b110010010110: bitmap = 51'b111111111111111000000000000000000000001111111111111;
        12'b110010010111: bitmap = 51'b111111111111110000000000000000000000011111111111111;
        12'b110010011000: bitmap = 51'b111111111111110000000000000000000000011111111111111;
        12'b110010011001: bitmap = 51'b111111111111100000000011111000000000111111111111111;
        12'b110010011010: bitmap = 51'b111111111111100000000111111100000000111111111111111;
        12'b110010011011: bitmap = 51'b111111111111000000001111111110000000011111111111111;
        12'b110010011100: bitmap = 51'b111111111111000000011111111111000000011111111111111;
        12'b110010011101: bitmap = 51'b111111111111000000011111111111000000011111111111111;
        12'b110010011110: bitmap = 51'b111111111111000000011111111111000000011111111111111;
        12'b110010011111: bitmap = 51'b111111111111000000011111111111000000011111111111111;
        12'b110010100000: bitmap = 51'b111111111111000000011111111111000000011111111111111;
        12'b110010100001: bitmap = 51'b111111111111000000001111111110000000011111111111111;
        12'b110010100010: bitmap = 51'b111111111111100000000111111100000000111111111111111;
        12'b110010100011: bitmap = 51'b111111111111100000000011111000000000111111111111111;
        12'b110010100100: bitmap = 51'b111111111111100000000000000000000001111111111111111;
        12'b110010100101: bitmap = 51'b111111111111110000000000000000000001111111111111111;
        12'b110010100110: bitmap = 51'b111111111111111000000000000000000011111111111111111;
        12'b110010100111: bitmap = 51'b111111111111111100000000000000000111111111111111111;
        12'b110010101000: bitmap = 51'b111111111111111110000000000000001111111111111111111;
        12'b110010101001: bitmap = 51'b111111111111111111100000000000111111111111111111111;
        12'b110010101010: bitmap = 51'b111111111111111111111000000011111111111111111111111;
        12'b110010101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110010101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110010101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b110010101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b110010101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b110010110000: bitmap = 51'b000001111111111111111111111111111111111111111000000;
        12'b110010110001: bitmap = 51'b000000011111111111111111111111111111111111100000000;
        12'b110010110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b110010110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b110010110100: bitmap = 51'b000000000000111111111111111111111111110000000000000;
        12'b110010110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b110010110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b110010110111: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b110010111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b110010111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b110010111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b110010111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        
        12'b110011000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b110011000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b110011000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b110011000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b110011000100: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b110011000101: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b110011000110: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b110011000111: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b110011001000: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b110011001001: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b110011001010: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b110011001011: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b110011001100: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b110011001101: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b110011001110: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b110011001111: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110011010000: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110011010001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110011010010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110011010011: bitmap = 51'b111111111111111111111100000001111111111111111111111;
        12'b110011010100: bitmap = 51'b111111111111111111110000000000011111111111111111111;
        12'b110011010101: bitmap = 51'b111111111111111111100000000000001111111111111111111;
        12'b110011010110: bitmap = 51'b111111111111111110000000000000000011111111111111111;
        12'b110011010111: bitmap = 51'b111111111111111110000000000000000000000000000000000;
        12'b110011011000: bitmap = 51'b111111111111101000000000000000000000000000000000000;
        12'b110011011001: bitmap = 51'b111111111111111000000001111000000000000000000000000;
        12'b110011011010: bitmap = 51'b111111111111111000000011111100000000000000000000000;
        12'b110011011011: bitmap = 51'b111111111111110000000111111110000000000000000000000;
        12'b110011011100: bitmap = 51'b111111111111110000001111111111000000000000000000000;
        12'b110011011101: bitmap = 51'b111111111111110000001111111111000000000000000000000;
        12'b110011011110: bitmap = 51'b111111111111110000001111111111000000000000000000000;
        12'b110011011111: bitmap = 51'b111111111111110000001111111111000000000000000000000;
        12'b110011100000: bitmap = 51'b111111111111110000000111111110000000000000000000000;
        12'b110011100001: bitmap = 51'b111111111111111000000011111100000000000000000000000;
        12'b110011100010: bitmap = 51'b111111111111111000000001111000000000000000000000000;
        12'b110011100011: bitmap = 51'b111111111111111100000000000000000000000000000000000;
        12'b110011100100: bitmap = 51'b111111111111111110000000000000000000000000000000000;
        12'b110011100101: bitmap = 51'b111111111111111110000000000000000011111111111111111;
        12'b110011100110: bitmap = 51'b111111111111111111100000000000001111111111111111111;
        12'b110011100111: bitmap = 51'b111111111111111111110000000000011111111111111111111;
        12'b110011101000: bitmap = 51'b111111111111111111111100000001111111111111111111111;
        12'b110011101001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110011101010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110011101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110011101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b110011101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b110011101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b110011101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b110011110000: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b110011110001: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b110011110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b110011110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b110011110100: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b110011110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b110011110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b110011110111: bitmap = 51'b000000000000000000111111111111111000000000000000000;
        12'b110011111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b110011111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b110011111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b110011111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        
      //shape 7 
        12'b111000000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b111000000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b111000000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b111000000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b111000000100: bitmap = 51'b000000000000000000011111111111110000000000000000000;
        12'b111000000101: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b111000000110: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b111000000111: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b111000001000: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b111000001001: bitmap = 51'b000000000000000000000011111110000000000000000000000;
        12'b111000001010: bitmap = 51'b000000000000000000000011111110000000000000000000000;
        12'b111000001011: bitmap = 51'b000000100000000000000001111100000000000000001000000;
        12'b111000001100: bitmap = 51'b000011110000000000000000111000000000000000011110000;
        12'b111000001101: bitmap = 51'b000111110000000000000000000000000000000000011111000;
        12'b111000001110: bitmap = 51'b011111111000000000000000000000000000000000111111110;
        12'b111000001111: bitmap = 51'b111111111000000000000000000000000000000000111111111;
        12'b111000010000: bitmap = 51'b111111111100000000000000000000000000000001111111111;
        12'b111000010001: bitmap = 51'b111111111100000000000000000000000000000001111111111;
        12'b111000010010: bitmap = 51'b111111111110000000000000000000000000000011111111111;
        12'b111000010011: bitmap = 51'b111111111111000000000000000000000000000111111111111;
        12'b111000010100: bitmap = 51'b111111111111000000000000000000000000000111111111111;
        12'b111000010101: bitmap = 51'b111111111111100000000000000000000000001111111111111;
        12'b111000010110: bitmap = 51'b111111111111100000000000000000000000001111111111111;
        12'b111000010111: bitmap = 51'b111111111111110000000000000000000000011111111111111;
        12'b111000011000: bitmap = 51'b111111111111110000000000000000000000011111111111111;
        12'b111000011001: bitmap = 51'b111111111111111000000000000000000000111111111111111;
        12'b111000011010: bitmap = 51'b111111111111111100000000000000000001111111111111111;
        12'b111000011011: bitmap = 51'b111111111111111100000000000000000001111111111111111;
        12'b111000011100: bitmap = 51'b111111111111111110000000000000000011111111111111111;
        12'b111000011101: bitmap = 51'b111111111111111110000000000000000011111111111111111;
        12'b111000011110: bitmap = 51'b111111111111111110000000000000000111111111111111111;
        12'b111000011111: bitmap = 51'b111111111111111110000000000000000111111111111111111;
        12'b111000100000: bitmap = 51'b111111111111111100000000000000001111111111111111111;
        12'b111000100001: bitmap = 51'b111111111111111100000000000000001111111111111111111;
        12'b111000100010: bitmap = 51'b111111111111111000000000000000011111111111111111111;
        12'b111000100011: bitmap = 51'b111111111111110000000000000000111111111111111111111;
        12'b111000100100: bitmap = 51'b111111111111110000000000000000111111111111111111111;
        12'b111000100101: bitmap = 51'b111111111111100000000000000001111111111111111111111;
        12'b111000100110: bitmap = 51'b111111111111100000000000000001111111111111111111111;
        12'b111000100111: bitmap = 51'b111111111111000000000000000011111111111111111111111;
        12'b111000101000: bitmap = 51'b111111111111000000000000000011111111111111111111111;
        12'b111000101001: bitmap = 51'b111111111110000000000000000111111111111111111111111;
        12'b111000101010: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b111000101011: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b111000101100: bitmap = 51'b111111111000000000000000011111111111111111111111111;
        12'b111000101101: bitmap = 51'b011111111000000000000000011111111111111111111111110;
        12'b111000101110: bitmap = 51'b000111110000000000000000111111111111111111111111000;
        12'b111000101111: bitmap = 51'b000011110000000000000000111111111111111111111110000;
        12'b111000110000: bitmap = 51'b000000100000000000000001111111111111111111111000000;
        12'b111000110001: bitmap = 51'b000000000000000000000011111111111111111111100000000;
        12'b111000110010: bitmap = 51'b000000000000000000000011111111111111111111000000000;
        12'b111000110011: bitmap = 51'b000000000000000000000111111111111111111100000000000;
        12'b111000110100: bitmap = 51'b000000000000000000000111111111111111110000000000000;
        12'b111000110101: bitmap = 51'b000000000000000000001111111111111111100000000000000;
        12'b111000110110: bitmap = 51'b000000000000000000001111111111111110000000000000000;
        12'b111000110111: bitmap = 51'b000000000000000000011111111111110000000000000000000;
        12'b111000111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b111000111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b111000111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b111000111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        
        
        12'b111001000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b111001000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b111001000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b111001000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b111001000100: bitmap = 51'b000000000000000000111111111111110000000000000000000;
        12'b111001000101: bitmap = 51'b000000000000000011111111111111100000000000000000000;
        12'b111001000110: bitmap = 51'b000000000000001111111111111111100000000000000000000;
        12'b111001000111: bitmap = 51'b000000000000011111111111111111000000000000000000000;
        12'b111001001000: bitmap = 51'b000000000001111111111111111111000000000000000000000;
        12'b111001001001: bitmap = 51'b000000000111111111111111111110000000000000000000000;
        12'b111001001010: bitmap = 51'b000000001111111111111111111110000000000000000000000;
        12'b111001001011: bitmap = 51'b000000111111111111111111111100000000000000001000000;
        12'b111001001100: bitmap = 51'b000011111111111111111111111000000000000000011110000;
        12'b111001001101: bitmap = 51'b000111111111111111111111111000000000000000011111000;
        12'b111001001110: bitmap = 51'b011111111111111111111111110000000000000000111111110;
        12'b111001001111: bitmap = 51'b111111111111111111111111110000000000000000111111111;
        12'b111001010000: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b111001010001: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b111001010010: bitmap = 51'b111111111111111111111111000000000000000011111111111;
        12'b111001010011: bitmap = 51'b111111111111111111111110000000000000000011111111111;
        12'b111001010100: bitmap = 51'b111111111111111111111110000000000000000011111111111;
        12'b111001010101: bitmap = 51'b111111111111111111111100000000000000000011111111111;
        12'b111001010110: bitmap = 51'b111111111111111111111100000000000000000001111111111;
        12'b111001010111: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111001011000: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111001011001: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111001011010: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111001011011: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111001011100: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111001011101: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111001011110: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111001011111: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111001100000: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111001100001: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111001100010: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111001100011: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111001100100: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111001100101: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b111001100110: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b111001100111: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b111001101000: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b111001101001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b111001101010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b111001101011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b111001101100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b111001101101: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b111001101110: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b111001101111: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b111001110000: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b111001110001: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b111001110010: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b111001110011: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b111001110100: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b111001110101: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b111001110110: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b111001110111: bitmap = 51'b000000000000000000011111111111111000000000000000000;
        12'b111001111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b111001111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b111001111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b111001111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        
        12'b111010000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b111010000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b111010000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b111010000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b111010000100: bitmap = 51'b000000000000000000011111111111111000000000000000000;
        12'b111010000101: bitmap = 51'b000000000000000000001111111111111110000000000000000;
        12'b111010000110: bitmap = 51'b000000000000000000001111111111111111100000000000000;
        12'b111010000111: bitmap = 51'b000000000000000000000111111111111111110000000000000;
        12'b111010001000: bitmap = 51'b000000000000000000000111111111111111111100000000000;
        12'b111010001001: bitmap = 51'b000000000000000000000011111111111111111111000000000;
        12'b111010001010: bitmap = 51'b000000000000000000000011111111111111111111100000000;
        12'b111010001011: bitmap = 51'b000000100000000000000001111111111111111111111000000;
        12'b111010001100: bitmap = 51'b000011110000000000000000111111111111111111111110000;
        12'b111010001101: bitmap = 51'b000111110000000000000000111111111111111111111111000;
        12'b111010001110: bitmap = 51'b011111111000000000000000011111111111111111111111110;
        12'b111010001111: bitmap = 51'b111111111000000000000000011111111111111111111111111;
        12'b111010010000: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b111010010001: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b111010010010: bitmap = 51'b111111111110000000000000000111111111111111111111111;
        12'b111010010011: bitmap = 51'b111111111111000000000000000011111111111111111111111;
        12'b111010010100: bitmap = 51'b111111111111000000000000000011111111111111111111111;
        12'b111010010101: bitmap = 51'b111111111111100000000000000001111111111111111111111;
        12'b111010010110: bitmap = 51'b111111111111100000000000000001111111111111111111111;
        12'b111010010111: bitmap = 51'b111111111111110000000000000000000000000000000000000;
        12'b111010011000: bitmap = 51'b111111111111110000000000000000000000000000000000000;
        12'b111010011001: bitmap = 51'b111111111111111000000000000000000000000000000000000;
        12'b111010011010: bitmap = 51'b111111111111111100000000000000000000000000000000000;
        12'b111010011011: bitmap = 51'b111111111111111100000000000000000000000000000000000;
        12'b111010011100: bitmap = 51'b111111111111111110000000000000000000000000000000000;
        12'b111010011101: bitmap = 51'b111111111111111110000000000000000000000000000000000;
        12'b111010011110: bitmap = 51'b111111111111111111000000000000000000000000000000000;
        12'b111010011111: bitmap = 51'b111111111111111111000000000000000000000000000000000;
        12'b111010100000: bitmap = 51'b111111111111111111100000000000000000000000000000000;
        12'b111010100001: bitmap = 51'b111111111111111111100000000000000000000000000000000;
        12'b111010100010: bitmap = 51'b111111111111111111110000000000000000000000000000000;
        12'b111010100011: bitmap = 51'b111111111111111111111000000000000000000000000000000;
        12'b111010100100: bitmap = 51'b111111111111111111111000000000000000000000000000000;
        12'b111010100101: bitmap = 51'b111111111111111111111100000000000000000001111111111;
        12'b111010100110: bitmap = 51'b111111111111111111111100000000000000000011111111111;
        12'b111010100111: bitmap = 51'b111111111111111111111110000000000000000011111111111;
        12'b111010101000: bitmap = 51'b111111111111111111111110000000000000000011111111111;
        12'b111010101001: bitmap = 51'b111111111111111111111111000000000000000011111111111;
        12'b111010101010: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b111010101011: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b111010101100: bitmap = 51'b111111111111111111111111110000000000000000111111111;
        12'b111010101101: bitmap = 51'b011111111111111111111111110000000000000000111111110;
        12'b111010101110: bitmap = 51'b000111111111111111111111111000000000000000011111000;
        12'b111010101111: bitmap = 51'b000011111111111111111111111000000000000000011110000;
        12'b111010110000: bitmap = 51'b000000111111111111111111111100000000000000001000000;
        12'b111010110001: bitmap = 51'b000000001111111111111111111110000000000000000000000;
        12'b111010110010: bitmap = 51'b000000000111111111111111111110000000000000000000000;
        12'b111010110011: bitmap = 51'b000000000001111111111111111111000000000000000000000;
        12'b111010110100: bitmap = 51'b000000000000011111111111111111000000000000000000000;
        12'b111010110101: bitmap = 51'b000000000000001111111111111111100000000000000000000;
        12'b111010110110: bitmap = 51'b000000000000000011111111111111100000000000000000000;
        12'b111010110111: bitmap = 51'b000000000000000000111111111111110000000000000000000;
        12'b111010111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b111010111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b111010111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b111010111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        
        12'b111011000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b111011000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b111011000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b111011000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b111011000100: bitmap = 51'b000000000000000000011111111111110000000000000000000;
        12'b111011000101: bitmap = 51'b000000000000000011111111111111100000000000000000000;
        12'b111011000110: bitmap = 51'b000000000000001111111111111111100000000000000000000;
        12'b111011000111: bitmap = 51'b000000000000011111111111111111000000000000000000000;
        12'b111011001000: bitmap = 51'b000000000001111111111111111111000000000000000000000;
        12'b111011001001: bitmap = 51'b000000000111111111111111111110000000000000000000000;
        12'b111011001010: bitmap = 51'b000000001111111111111111111110000000000000000000000;
        12'b111011001011: bitmap = 51'b000000111111111111111111111100000000000000001000000;
        12'b111011001100: bitmap = 51'b000011111111111111111111111000000000000000011110000;
        12'b111011001101: bitmap = 51'b000111111111111111111111111000000000000000011111000;
        12'b111011001110: bitmap = 51'b011111111111111111111111110000000000000000111111110;
        12'b111011001111: bitmap = 51'b111111111111111111111111110000000000000000111111111;
        12'b111011010000: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b111011010001: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b111011010010: bitmap = 51'b111111111111111111111111000000000000000011111111111;
        12'b111011010011: bitmap = 51'b111111111111111111111110000000000000000111111111111;
        12'b111011010100: bitmap = 51'b111111111111111111111110000000000000000111111111111;
        12'b111011010101: bitmap = 51'b111111111111111111111100000000000000001111111111111;
        12'b111011010110: bitmap = 51'b111111111111111111111100000000000000001111111111111;
        12'b111011010111: bitmap = 51'b111111111111111111111000000000000000011111111111111;
        12'b111011011000: bitmap = 51'b111111111111111111111000000000000000011111111111111;
        12'b111011011001: bitmap = 51'b111111111111111111110000000000000000111111111111111;
        12'b111011011010: bitmap = 51'b111111111111111111100000000000000001111111111111111;
        12'b111011011011: bitmap = 51'b111111111111111111100000000000000001111111111111111;
        12'b111011011100: bitmap = 51'b111111111111111111000000000000000011111111111111111;
        12'b111011011101: bitmap = 51'b111111111111111111000000000000000011111111111111111;
        12'b111011011110: bitmap = 51'b111111111111111110000000000000000011111111111111111;
        12'b111011011111: bitmap = 51'b111111111111111110000000000000000011111111111111111;
        12'b111011100000: bitmap = 51'b111111111111111100000000000000000001111111111111111;
        12'b111011100001: bitmap = 51'b111111111111111100000000000000000001111111111111111;
        12'b111011100010: bitmap = 51'b111111111111111000000000000000000000111111111111111;
        12'b111011100011: bitmap = 51'b111111111111110000000000000000000000011111111111111;
        12'b111011100100: bitmap = 51'b111111111111110000000000000000000000011111111111111;
        12'b111011100101: bitmap = 51'b111111111111100000000000000000000000001111111111111;
        12'b111011100110: bitmap = 51'b111111111111100000000000000000000000001111111111111;
        12'b111011100111: bitmap = 51'b111111111111000000000000000000000000000111111111111;
        12'b111011101000: bitmap = 51'b111111111111000000000000000000000000000111111111111;
        12'b111011101001: bitmap = 51'b111111111110000000000000000000000000000011111111111;
        12'b111011101010: bitmap = 51'b111111111100000000000000000000000000000001111111111;
        12'b111011101011: bitmap = 51'b111111111100000000000000000000000000000001111111111;
        12'b111011101100: bitmap = 51'b111111111000000000000000000000000000000000111111111;
        12'b111011101101: bitmap = 51'b011111111000000000000000000000000000000000111111110;
        12'b111011101110: bitmap = 51'b000111110000000000000000000000000000000000011111000;
        12'b111011101111: bitmap = 51'b000011110000000000000000111000000000000000011110000;
        12'b111011110000: bitmap = 51'b000000100000000000000001111100000000000000001000000;
        12'b111011110001: bitmap = 51'b000000000000000000000011111110000000000000000000000;
        12'b111011110010: bitmap = 51'b000000000000000000000011111110000000000000000000000;
        12'b111011110011: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b111011110100: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b111011110101: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b111011110110: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b111011110111: bitmap = 51'b000000000000000000011111111111110000000000000000000;
        12'b111011111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b111011111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b111011111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b111011111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;

        12'b111100000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b111100000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b111100000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b111100000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b111100000100: bitmap = 51'b000000000000000000111111111111110000000000000000000;
        12'b111100000101: bitmap = 51'b000000000000000011111111111111111110000000000000000;
        12'b111100000110: bitmap = 51'b000000000000001111111111111111111111100000000000000;
        12'b111100000111: bitmap = 51'b000000000000011111111111111111111111110000000000000;
        12'b111100001000: bitmap = 51'b000000000001111111111111111111111111111100000000000;
        12'b111100001001: bitmap = 51'b000000000111111111111111111111111111111111000000000;
        12'b111100001010: bitmap = 51'b000000001111111111111111111111111111111111100000000;
        12'b111100001011: bitmap = 51'b000000111111111111111111111111111111111111111000000;
        12'b111100001100: bitmap = 51'b000011111111111111111111111111111111111111111110000;
        12'b111100001101: bitmap = 51'b000111111111111111111111111111111111111111111111000;
        12'b111100001110: bitmap = 51'b011111111111111111111111111111111111111111111111110;
        12'b111100001111: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b111100010000: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b111100010001: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b111100010010: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b111100010011: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b111100010100: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b111100010101: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b111100010110: bitmap = 51'b111111111111111111111111111111111111111111111111111;
        12'b111100010111: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111100011000: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111100011001: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111100011010: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111100011011: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111100011100: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111100011101: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111100011110: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111100011111: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111100100000: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111100100001: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111100100010: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111100100011: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111100100100: bitmap = 51'b000000000000000000000000000000000000000000000000000;
        12'b111100100101: bitmap = 51'b111111111100000000000000000001111111111111111111111;
        12'b111100100110: bitmap = 51'b111111111110000000000000000001111111111111111111111;
        12'b111100100111: bitmap = 51'b111111111110000000000000000011111111111111111111111;
        12'b111100101000: bitmap = 51'b111111111110000000000000000011111111111111111111111;
        12'b111100101001: bitmap = 51'b111111111110000000000000000111111111111111111111111;
        12'b111100101010: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b111100101011: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b111100101100: bitmap = 51'b111111111000000000000000011111111111111111111111111;
        12'b111100101101: bitmap = 51'b011111111000000000000000011111111111111111111111110;
        12'b111100101110: bitmap = 51'b000111110000000000000000111111111111111111111111000;
        12'b111100101111: bitmap = 51'b000011110000000000000000111111111111111111111110000;
        12'b111100110000: bitmap = 51'b000000100000000000000001111111111111111111111000000;
        12'b111100110001: bitmap = 51'b000000000000000000000011111111111111111111100000000;
        12'b111100110010: bitmap = 51'b000000000000000000000011111111111111111111000000000;
        12'b111100110011: bitmap = 51'b000000000000000000000111111111111111111100000000000;
        12'b111100110100: bitmap = 51'b000000000000000000000111111111111111110000000000000;
        12'b111100110101: bitmap = 51'b000000000000000000001111111111111111100000000000000;
        12'b111100110110: bitmap = 51'b000000000000000000001111111111111110000000000000000;
        12'b111100110111: bitmap = 51'b000000000000000000011111111111111000000000000000000;
        12'b111100111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b111100111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b111100111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b111100111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;

        12'b111101000000: bitmap = 51'b000000000000000000000000010000000000000000000000000;
        12'b111101000001: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b111101000010: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b111101000011: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b111101000100: bitmap = 51'b000000000000000000011111111111111000000000000000000;
        12'b111101000101: bitmap = 51'b000000000000000000001111111111111110000000000000000;
        12'b111101000110: bitmap = 51'b000000000000000000001111111111111111100000000000000;
        12'b111101000111: bitmap = 51'b000000000000000000000111111111111111110000000000000;
        12'b111101001000: bitmap = 51'b000000000000000000000111111111111111111100000000000;
        12'b111101001001: bitmap = 51'b000000000000000000000011111111111111111111000000000;
        12'b111101001010: bitmap = 51'b000000000000000000000011111111111111111111100000000;
        12'b111101001011: bitmap = 51'b000000100000000000000001111111111111111111111000000;
        12'b111101001100: bitmap = 51'b000011110000000000000000111111111111111111111110000;
        12'b111101001101: bitmap = 51'b000111110000000000000000111111111111111111111111000;
        12'b111101001110: bitmap = 51'b011111111000000000000000011111111111111111111111110;
        12'b111101001111: bitmap = 51'b111111111000000000000000011111111111111111111111111;
        12'b111101010000: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b111101010001: bitmap = 51'b111111111100000000000000001111111111111111111111111;
        12'b111101010010: bitmap = 51'b111111111110000000000000000111111111111111111111111;
        12'b111101010011: bitmap = 51'b111111111110000000000000000011111111111111111111111;
        12'b111101010100: bitmap = 51'b111111111110000000000000000011111111111111111111111;
        12'b111101010101: bitmap = 51'b111111111110000000000000000001111111111111111111111;
        12'b111101010110: bitmap = 51'b111111111100000000000000000001111111111111111111111;
        12'b111101010111: bitmap = 51'b000000000000000000000000000000111111111111111111111;
        12'b111101011000: bitmap = 51'b000000000000000000000000000000111111111111111111111;
        12'b111101011001: bitmap = 51'b000000000000000000000000000000011111111111111111111;
        12'b111101011010: bitmap = 51'b000000000000000000000000000000001111111111111111111;
        12'b111101011011: bitmap = 51'b000000000000000000000000000000001111111111111111111;
        12'b111101011100: bitmap = 51'b000000000000000000000000000000000111111111111111111;
        12'b111101011101: bitmap = 51'b000000000000000000000000000000000111111111111111111;
        12'b111101011110: bitmap = 51'b000000000000000000000000000000000011111111111111111;
        12'b111101011111: bitmap = 51'b000000000000000000000000000000000011111111111111111;
        12'b111101100000: bitmap = 51'b000000000000000000000000000000000001111111111111111;
        12'b111101100001: bitmap = 51'b000000000000000000000000000000000001111111111111111;
        12'b111101100010: bitmap = 51'b000000000000000000000000000000000000111111111111111;
        12'b111101100011: bitmap = 51'b000000000000000000000000000000000000011111111111111;
        12'b111101100100: bitmap = 51'b000000000000000000000000000000000000011111111111111;
        12'b111101100101: bitmap = 51'b111111111111111111111100000000000000001111111111111;
        12'b111101100110: bitmap = 51'b111111111111111111111100000000000000001111111111111;
        12'b111101100111: bitmap = 51'b111111111111111111111110000000000000000111111111111;
        12'b111101101000: bitmap = 51'b111111111111111111111110000000000000000111111111111;
        12'b111101101001: bitmap = 51'b111111111111111111111111000000000000000011111111111;
        12'b111101101010: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b111101101011: bitmap = 51'b111111111111111111111111100000000000000001111111111;
        12'b111101101100: bitmap = 51'b111111111111111111111111110000000000000000111111111;
        12'b111101101101: bitmap = 51'b011111111111111111111111110000000000000000111111110;
        12'b111101101110: bitmap = 51'b000111111111111111111111111000000000000000011111000;
        12'b111101101111: bitmap = 51'b000011111111111111111111111000000000000000011110000;
        12'b111101110000: bitmap = 51'b000000111111111111111111111100000000000000001000000;
        12'b111101110001: bitmap = 51'b000000001111111111111111111110000000000000000000000;
        12'b111101110010: bitmap = 51'b000000000111111111111111111110000000000000000000000;
        12'b111101110011: bitmap = 51'b000000000001111111111111111111000000000000000000000;
        12'b111101110100: bitmap = 51'b000000000000011111111111111111000000000000000000000;
        12'b111101110101: bitmap = 51'b000000000000001111111111111111100000000000000000000;
        12'b111101110110: bitmap = 51'b000000000000000011111111111111100000000000000000000;
        12'b111101110111: bitmap = 51'b000000000000000000111111111111110000000000000000000;
        12'b111101111000: bitmap = 51'b000000000000000000001111111111100000000000000000000;
        12'b111101111001: bitmap = 51'b000000000000000000000111111111000000000000000000000;
        12'b111101111010: bitmap = 51'b000000000000000000000001111100000000000000000000000;
        12'b111101111011: bitmap = 51'b000000000000000000000000010000000000000000000000000;
    endcase
  end
  
endmodule