module shape5base (
    input wire clk,  // clock
    input [2:0] orientation,
    input wire[5:0] address,
    output reg [50:0] outdata
  );
  
  (* rom_style = "block" *)
  
  reg [5:0] address_reg;
  reg[2:0] orientreg;
  
  always @(posedge clk) begin
    address_reg <= address;
    orientreg <= orientation;
    
  end

  /* Combinational Logic */
  always @* begin
      case({orientreg,address_reg})
          9'b000000000: outdata = 51'b000000000000000000000000010000000000000000000000000;
          9'b000000001: outdata = 51'b000000000000000000000001111100000000000000000000000;
          9'b000000010: outdata = 51'b000000000000000000000111111111000000000000000000000;
          9'b000000011: outdata = 51'b000000000000000000001111111111100000000000000000000;
          9'b000000100: outdata = 51'b000000000000000000111111111111111000000000000000000;
          9'b000000101: outdata = 51'b000000000000000011111111111111111110000000000000000;
          9'b000000110: outdata = 51'b000000000000001111111111111111111111100000000000000;
          9'b000000111: outdata = 51'b000000000000011111111111111111111111110000000000000;
          9'b000001000: outdata = 51'b000000000001111111111111111111111111111100000000000;
          9'b000001001: outdata = 51'b000000000111111111111111111111111111111111000000000;
          9'b000001010: outdata = 51'b000000001111111111111111111111111111111111100000000;
          9'b000001011: outdata = 51'b000000111111111111111111111111111111111111111000000;
          9'b000001100: outdata = 51'b000011111111111111111111111111111111111111111110000;
          9'b000001101: outdata = 51'b000111111111111111111111111111111111111111111111000;
          9'b000001110: outdata = 51'b011111111111111111111111111111111111111111111111110;
          9'b000001111: outdata = 51'b111111111111111111111111111111111111111111111111111;
          9'b000010000: outdata = 51'b111111111111111111111111111111111111111111111111111;
          9'b000010001: outdata = 51'b111111111111111111111111111111111111111111111111111;
          9'b000010010: outdata = 51'b111111111111111111111111111111111111111111111111111;
          9'b000010011: outdata = 51'b111111111111111111111100000001111111111111111111111;
          9'b000010100: outdata = 51'b111111111111111111110000000000011111111111111111111;
          9'b000010101: outdata = 51'b111111111111111111100000000000001111111111111111111;
          9'b000010110: outdata = 51'b111111111111111110000000000000000011111111111111111;
          9'b000010111: outdata = 51'b000000000000000000000000000000000011111111111111111;
          9'b000011000: outdata = 51'b000000000000000000000000000000000000101111111111111;
          9'b000011001: outdata = 51'b000000000000000000000000000000000000111111111111111;
          9'b000011010: outdata = 51'b000000000000000000000000000000000000111111111111111;
          9'b000011011: outdata = 51'b000000000000000000000000000000000000011111111111111;
          9'b000011100: outdata = 51'b000000000000000000000000000000000000011111111111111;
          9'b000011101: outdata = 51'b000000000000000000000000000000000000011111111111111;
          9'b000011110: outdata = 51'b000000000000000000000000000000000000011111111111111;
          9'b000011111: outdata = 51'b000000000000000000000000000000000000011111111111111;
          9'b000100000: outdata = 51'b000000000000000000000000000000000000011111111111111;
          9'b000100001: outdata = 51'b000000000000000000000000000000000000111111111111111;
          9'b000100010: outdata = 51'b000000000000000000000000000000000000111111111111111;
          9'b000100011: outdata = 51'b000000000000000000000000000000000001111111111111111;
          9'b000100100: outdata = 51'b000000000000000000000000000000000011111111111111111;
          9'b000100101: outdata = 51'b111111111111111110000000000000000011111111111111111;
          9'b000100110: outdata = 51'b111111111111111111100000000000001111111111111111111;
          9'b000100111: outdata = 51'b111111111111111111110000000000011111111111111111111;
          9'b000101000: outdata = 51'b111111111111111111111100000001111111111111111111111;
          9'b000101001: outdata = 51'b111111111111111111111111111111111111111111111111111;
          9'b000101010: outdata = 51'b111111111111111111111111111111111111111111111111111;
          9'b000101011: outdata = 51'b111111111111111111111111111111111111111111111111111;
          9'b000101100: outdata = 51'b111111111111111111111111111111111111111111111111111;
          9'b000101101: outdata = 51'b011111111111111111111111111111111111111111111111110;
          9'b000101110: outdata = 51'b000111111111111111111111111111111111111111111111000;
          9'b000101111: outdata = 51'b000011111111111111111111111111111111111111111110000;
          9'b000110000: outdata = 51'b000000111111111111111111111111111111111111111000000;
          9'b000110001: outdata = 51'b000000001111111111111111111111111111111111100000000;
          9'b000110010: outdata = 51'b000000000111111111111111111111111111111111000000000;
          9'b000110011: outdata = 51'b000000000001111111111111111111111111111100000000000;
          9'b000110100: outdata = 51'b000000000000011111111111111111111111110000000000000;
          9'b000110101: outdata = 51'b000000000000001111111111111111111111100000000000000;
          9'b000110110: outdata = 51'b000000000000000011111111111111111110000000000000000;
          9'b000110111: outdata = 51'b000000000000000000111111111111111000000000000000000;
          9'b000111000: outdata = 51'b000000000000000000001111111111100000000000000000000;
          9'b000111001: outdata = 51'b000000000000000000000111111111000000000000000000000;
          9'b000111010: outdata = 51'b000000000000000000000001111100000000000000000000000;
          9'b000111011: outdata = 51'b000000000000000000000000010000000000000000000000000;
          
          
          
          9'b001000000: outdata = 51'b000000000000000000000000010000000000000000000000000;
          9'b001000001: outdata = 51'b000000000000000000000001111100000000000000000000000;
          9'b001000010: outdata = 51'b000000000000000000000111111111000000000000000000000;
          9'b001000011: outdata = 51'b000000000000000000001111111111100000000000000000000;
          9'b001000100: outdata = 51'b000000000000000000011111111111111000000000000000000;
          9'b001000101: outdata = 51'b000000000000000000001111111111111110000000000000000;
          9'b001000110: outdata = 51'b000000000000000000001111111111111111100000000000000;
          9'b001000111: outdata = 51'b000000000000000000000111111111111111110000000000000;
          9'b001001000: outdata = 51'b000000000000000000000111111111111111111100000000000;
          9'b001001001: outdata = 51'b000000000000000000000011111111111111111111000000000;
          9'b001001010: outdata = 51'b000000000000000000000011111111111111111111100000000;
          9'b001001011: outdata = 51'b000000100000000000000001111111111111111111111000000;
          9'b001001100: outdata = 51'b000011110000000000000000111111111111111111111110000;
          9'b001001101: outdata = 51'b000111110000000000000000111111111111111111111111000;
          9'b001001110: outdata = 51'b011111111000000000000000011111111111111111111111110;
          9'b001001111: outdata = 51'b111111111000000000000000011111111111111111111111111;
          9'b001010000: outdata = 51'b111111111100000000000000001111111111111111111111111;
          9'b001010001: outdata = 51'b111111111100000000000000000111111111111111111111111;
          9'b001010010: outdata = 51'b111111111110000000000000000011111111111111111111111;
          9'b001010011: outdata = 51'b111111111110000000000000000000001111111111111111111;
          9'b001010100: outdata = 51'b111111111111000000000000000000000011111111111111111;
          9'b001010101: outdata = 51'b111111111111100000000000000000000001111111111111111;
          9'b001010110: outdata = 51'b111111111111100000000000000000000000111111111111111;
          9'b001010111: outdata = 51'b111111111111110000000000000000000000011111111111111;
          9'b001011000: outdata = 51'b111111111111110000000000000000000000011111111111111;
          9'b001011001: outdata = 51'b111111111111111000000000000000000000001111111111111;
          9'b001011010: outdata = 51'b111111111111111000000000000000000000001111111111111;
          9'b001011011: outdata = 51'b111111111111111000000000000000000000000111111111111;
          9'b001011100: outdata = 51'b111111111111110000000000000000000000000111111111111;
          9'b001011101: outdata = 51'b111111111111110000000000000000000000000111111111111;
          9'b001011110: outdata = 51'b111111111111110000000000000000000000000111111111111;
          9'b001011111: outdata = 51'b111111111111110000000000000000000000000111111111111;
          9'b001100000: outdata = 51'b111111111111110000000000000000000000000111111111111;
          9'b001100001: outdata = 51'b111111111111110000000000000000000000000111111111111;
          9'b001100010: outdata = 51'b111111111111111000000000000000000000001111111111111;
          9'b001100011: outdata = 51'b111111111111111000000000000000000000001111111111111;
          9'b001100100: outdata = 51'b111111111111111100000000000000000000001111111111111;
          9'b001100101: outdata = 51'b111111111111111100000000000000000000011111111111111;
          9'b001100110: outdata = 51'b111111111111111110000000000000000000111111111111111;
          9'b001100111: outdata = 51'b111111111111111111000000000000000001111111111111111;
          9'b001101000: outdata = 51'b111111111111111111100000000000000011111111111111111;
          9'b001101001: outdata = 51'b111111111111111111111000000000001111111111111111111;
          9'b001101010: outdata = 51'b111111111111111111111110000000111111111111111111111;
          9'b001101011: outdata = 51'b111111111111111111111111111111111111111111111111111;
          9'b001101100: outdata = 51'b111111111111111111111111111111111111111111111111111;
          9'b001101101: outdata = 51'b011111111111111111111111111111111111111111111111110;
          9'b001101110: outdata = 51'b000111111111111111111111111111111111111111111111000;
          9'b001101111: outdata = 51'b000011111111111111111111111111111111111111111110000;
          9'b001110000: outdata = 51'b000000111111111111111111111111111111111111111100000;
          9'b001110001: outdata = 51'b000000001111111111111111111111111111111111110000000;
          9'b001110010: outdata = 51'b000000000111111111111111111111111111111111000000000;
          9'b001110011: outdata = 51'b000000000001111111111111111111111111111100000000000;
          9'b001110100: outdata = 51'b000000000000011111111111111111111111111000000000000;
          9'b001110101: outdata = 51'b000000000000001111111111111111111111100000000000000;
          9'b001110110: outdata = 51'b000000000000000011111111111111111110000000000000000;
          9'b001110111: outdata = 51'b000000000000000000111111111111111000000000000000000;
          9'b001111000: outdata = 51'b000000000000000000001111111111100000000000000000000;
          9'b001111001: outdata = 51'b000000000000000000000111111111000000000000000000000;
          9'b001111010: outdata = 51'b000000000000000000000001111100000000000000000000000;
          9'b001111011: outdata = 51'b000000000000000000000000010000000000000000000000000;
          
          9'b011000000: outdata = 51'b000000000000000000000000010000000000000000000000000;
          9'b011000001: outdata = 51'b000000000000000000000001111100000000000000000000000;
          9'b011000010: outdata = 51'b000000000000000000000111111111000000000000000000000;
          9'b011000011: outdata = 51'b000000000000000000001111111111100000000000000000000;
          9'b011000100: outdata = 51'b000000000000000000111111111111110000000000000000000;
          9'b011000101: outdata = 51'b000000000000000011111111111111100000000000000000000;
          9'b011000110: outdata = 51'b000000000000001111111111111111100000000000000000000;
          9'b011000111: outdata = 51'b000000000000011111111111111111000000000000000000000;
          9'b011001000: outdata = 51'b000000000001111111111111111111000000000000000000000;
          9'b011001001: outdata = 51'b000000000111111111111111111110000000000000000000000;
          9'b011001010: outdata = 51'b000000001111111111111111111110000000000000000000000;
          9'b011001011: outdata = 51'b000000111111111111111111111100000000000000001000000;
          9'b011001100: outdata = 51'b000011111111111111111111111000000000000000011110000;
          9'b011001101: outdata = 51'b000111111111111111111111111000000000000000011111000;
          9'b011001110: outdata = 51'b011111111111111111111111110000000000000000111111110;
          9'b011001111: outdata = 51'b111111111111111111111111110000000000000000111111111;
          9'b011010000: outdata = 51'b111111111111111111111111100000000000000001111111111;
          9'b011010001: outdata = 51'b111111111111111111111111000000000000000001111111111;
          9'b011010010: outdata = 51'b111111111111111111111110000000000000000011111111111;
          9'b011010011: outdata = 51'b111111111111111111100000000000000000000011111111111;
          9'b011010100: outdata = 51'b111111111111111110000000000000000000000111111111111;
          9'b011010101: outdata = 51'b111111111111111100000000000000000000001111111111111;
          9'b011010110: outdata = 51'b111111111111111000000000000000000000001111111111111;
          9'b011010111: outdata = 51'b111111111111110000000000000000000000011111111111111;
          9'b011011000: outdata = 51'b111111111111110000000000000000000000011111111111111;
          9'b011011001: outdata = 51'b111111111111100000000000000000000000111111111111111;
          9'b011011010: outdata = 51'b111111111111100000000000000000000000111111111111111;
          9'b011011011: outdata = 51'b111111111111000000000000000000000000111111111111111;
          9'b011011100: outdata = 51'b111111111111000000000000000000000000011111111111111;
          9'b011011101: outdata = 51'b111111111111000000000000000000000000011111111111111;
          9'b011011110: outdata = 51'b111111111111000000000000000000000000011111111111111;
          9'b011011111: outdata = 51'b111111111111000000000000000000000000011111111111111;
          9'b011100000: outdata = 51'b111111111111000000000000000000000000011111111111111;
          9'b011100001: outdata = 51'b111111111111000000000000000000000000011111111111111;
          9'b011100010: outdata = 51'b111111111111100000000000000000000000111111111111111;
          9'b011100011: outdata = 51'b111111111111100000000000000000000000111111111111111;
          9'b011100100: outdata = 51'b111111111111100000000000000000000001111111111111111;
          9'b011100101: outdata = 51'b111111111111110000000000000000000001111111111111111;
          9'b011100110: outdata = 51'b111111111111111000000000000000000011111111111111111;
          9'b011100111: outdata = 51'b111111111111111100000000000000000111111111111111111;
          9'b011101000: outdata = 51'b111111111111111110000000000000001111111111111111111;
          9'b011101001: outdata = 51'b111111111111111111100000000000111111111111111111111;
          9'b011101010: outdata = 51'b111111111111111111111000000011111111111111111111111;
          9'b011101011: outdata = 51'b111111111111111111111111111111111111111111111111111;
          9'b011101100: outdata = 51'b111111111111111111111111111111111111111111111111111;
          9'b011101101: outdata = 51'b011111111111111111111111111111111111111111111111110;
          9'b011101110: outdata = 51'b000111111111111111111111111111111111111111111111000;
          9'b011101111: outdata = 51'b000011111111111111111111111111111111111111111110000;
          9'b011110000: outdata = 51'b000001111111111111111111111111111111111111111000000;
          9'b011110001: outdata = 51'b000000011111111111111111111111111111111111100000000;
          9'b011110010: outdata = 51'b000000000111111111111111111111111111111111000000000;
          9'b011110011: outdata = 51'b000000000001111111111111111111111111111100000000000;
          9'b011110100: outdata = 51'b000000000000111111111111111111111111110000000000000;
          9'b011110101: outdata = 51'b000000000000001111111111111111111111100000000000000;
          9'b011110110: outdata = 51'b000000000000000011111111111111111110000000000000000;
          9'b011110111: outdata = 51'b000000000000000000111111111111111000000000000000000;
          9'b011111000: outdata = 51'b000000000000000000001111111111100000000000000000000;
          9'b011111001: outdata = 51'b000000000000000000000111111111000000000000000000000;
          9'b011111010: outdata = 51'b000000000000000000000001111100000000000000000000000;
          9'b011111011: outdata = 51'b000000000000000000000000010000000000000000000000000;
          
          0: outdata = 51'b000000000000000000000000010000000000000000000000000;
          1: outdata = 51'b000000000000000000000001111100000000000000000000000;
          2: outdata = 51'b000000000000000000000111111111000000000000000000000;
          3: outdata = 51'b000000000000000000001111111111100000000000000000000;
          4: outdata = 51'b000000000000000000111111111111111000000000000000000;
          5: outdata = 51'b000000000000000011111111111111111110000000000000000;
          6: outdata = 51'b000000000000001111111111111111111111100000000000000;
          7: outdata = 51'b000000000000011111111111111111111111110000000000000;
          8: outdata = 51'b000000000001111111111111111111111111111100000000000;
          9: outdata = 51'b000000000111111111111111111111111111111111000000000;
          10: outdata = 51'b000000001111111111111111111111111111111111100000000;
          11: outdata = 51'b000000111111111111111111111111111111111111111000000;
          12: outdata = 51'b000011111111111111111111111111111111111111111110000;
          13: outdata = 51'b000111111111111111111111111111111111111111111111000;
          14: outdata = 51'b011111111111111111111111111111111111111111111111110;
          15: outdata = 51'b111111111111111111111111111111111111111111111111111;
          16: outdata = 51'b111111111111111111111111111111111111111111111111111;
          17: outdata = 51'b111111111111111111111111111111111111111111111111111;
          18: outdata = 51'b111111111111111111111111111111111111111111111111111;
          19: outdata = 51'b111111111111111111111100000001111111111111111111111;
          20: outdata = 51'b111111111111111111110000000000011111111111111111111;
          21: outdata = 51'b111111111111111111100000000000001111111111111111111;
          22: outdata = 51'b111111111111111110000000000000000011111111111111111;
          23: outdata = 51'b111111111111111110000000000000000000000000000000000;
          24: outdata = 51'b111111111111101000000000000000000000000000000000000;
          25: outdata = 51'b111111111111111000000000000000000000000000000000000;
          26: outdata = 51'b111111111111111000000000000000000000000000000000000;
          27: outdata = 51'b111111111111110000000000000000000000000000000000000;
          28: outdata = 51'b111111111111110000000000000000000000000000000000000;
          29: outdata = 51'b111111111111110000000000000000000000000000000000000;
          30: outdata = 51'b111111111111110000000000000000000000000000000000000;
          31: outdata = 51'b111111111111110000000000000000000000000000000000000;
          32: outdata = 51'b111111111111110000000000000000000000000000000000000;
          33: outdata = 51'b111111111111111000000000000000000000000000000000000;
          34: outdata = 51'b111111111111111000000000000000000000000000000000000;
          35: outdata = 51'b111111111111111100000000000000000000000000000000000;
          36: outdata = 51'b111111111111111110000000000000000000000000000000000;
          37: outdata = 51'b111111111111111110000000000000000011111111111111111;
          38: outdata = 51'b111111111111111111100000000000001111111111111111111;
          39: outdata = 51'b111111111111111111110000000000011111111111111111111;
          40: outdata = 51'b111111111111111111111100000001111111111111111111111;
          41: outdata = 51'b111111111111111111111111111111111111111111111111111;
          42: outdata = 51'b111111111111111111111111111111111111111111111111111;
          43: outdata = 51'b111111111111111111111111111111111111111111111111111;
          44: outdata = 51'b111111111111111111111111111111111111111111111111111;
          45: outdata = 51'b011111111111111111111111111111111111111111111111110;
          46: outdata = 51'b000111111111111111111111111111111111111111111111000;
          47: outdata = 51'b000011111111111111111111111111111111111111111110000;
          48: outdata = 51'b000000111111111111111111111111111111111111111000000;
          49: outdata = 51'b000000001111111111111111111111111111111111100000000;
          50: outdata = 51'b000000000111111111111111111111111111111111000000000;
          51: outdata = 51'b000000000001111111111111111111111111111100000000000;
          52: outdata = 51'b000000000000011111111111111111111111110000000000000;
          53: outdata = 51'b000000000000001111111111111111111111100000000000000;
          54: outdata = 51'b000000000000000011111111111111111110000000000000000;
          55: outdata = 51'b000000000000000000111111111111111000000000000000000;
          56: outdata = 51'b000000000000000000001111111111100000000000000000000;
          57: outdata = 51'b000000000000000000000111111111000000000000000000000;
          58: outdata = 51'b000000000000000000000001111100000000000000000000000;
          59: outdata = 51'b000000000000000000000000010000000000000000000000000;


          default: outdata = 0;
          
          endcase
  end
  
endmodule