module header (clk, en, address, bitmap); 
    input  clk;
    input   en;
    input wire[6:0] address;
    output reg [589:0] bitmap;
    reg [6:0]address_reg;
    
 always @(posedge clk)
 begin
   if (en)
     address_reg <= address;
 end

 always @(address_reg) 
 begin
    if (en)
       case(address_reg)
        0: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        1: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        2: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        3: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        4: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        6: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        7: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        8: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        9: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000;
        10: bitmap <= 590'b00000000000000000000000000100000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000010000000001000100000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000100000000000001000100000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000;
        11: bitmap <= 590'b00000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000100000001000000000000000100000000000000000000000001000000000000000000010000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000001010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000010001000000000000000000;
        12: bitmap <= 590'b10000000000100000000000000000000000000000000000000000000100010000000000000010000001000000000000000010010000000000000000010000000000000000001000000100000000000000001001000000000000000000000100000000000000010001000000000000000000010000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000001000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000001010000000000100;
        13: bitmap <= 590'b00000000000000000000000000000000010000010000000010100100000000000000000001000000000000000000000001001000000000000100000000000000000000000100000000000000000000000000100000000000010101000000000000000000000000000000000000000000000000000000000101010000000000000000000001001000000000000000000001000001000000001001000000000000000000000010100000000000000000000010100000000000100000000000000000000000001000000000000000000000000000010000000010010100000000000000000000100000010000000000000000100100000000001010000000000000000000000001000000000000000000000000000000000000100000000000000000000000010000;
        14: bitmap <= 590'b00000000001000000000000000000000000100000000000100000000000000000000100000010000000000000000000000000000001000001000100000000000000000000010000000000000000000000100000010000000000000100000000000000000010000000000000000000000010000100010000000000000000000000000000000100000000000000000000000010000100000000100100000000000000000000100000000000000000000000000000010000000010000100000000000001000000010000000000000000000010110000010000001000000000000000000100000000000001000000000000000010000101000000000100000000000000010000100000000000000000000000110000000100000010000000000000000001000001000;
        15: bitmap <= 590'b00110100000101000000000010000101000001000100000010010100000100100000010000001010000000101000000010000000000001000100110000010001000110000001000000000101010000010010000001000110000000010000010100100000000100000000010101000000001000000000000100001001000010110001010000011000000001010100010001000100010001000000010000000011001010000000100000000001010001011001000001000100000010010000100100000000001001000000010010000010000001000000001000000000000100010100010001010100000001010100000100010000000000001000010000010001010001000010101000000101010001000010010000000100000100010000100000000100000010;
        16: bitmap <= 590'b10010010010101000000001000000000011001000010001000000000000010010101001001001000000000001010001010100100000000100000001000000100010010000001011000000000100001000000010000000011000000000000000000010000000101000000000010100100001001001000000000100000000000001010001000000100000000000010000100000000000000101001001010001000100010000000010000000001000000000000100000000010101000001000100101000010001000100000000000100001001001001000000010101010000010100010000000001010000000100000001010001100000001000010001000010100001000000010100000000000100001000000010010000010000100001000010110100000000101;
        17: bitmap <= 590'b01000000000010101001100101000010100000010000000001010000000000000010000000100001000101010000000000001001000100000100000000000001000001000010000000000010000000010101000000000100001100000000010100100000010001000001010100000010100110010001011001000100000000100100000000100011000001010000010000010100000101000001000000000000011000000110100100011100010000010100110000010101000000000000000000110100010100011000101010000010100000010001111000010000000000010010001000010100000100010100010001000001000101010001010000000000000101100100010010001100000000010101000000010001001001000000000000010000010000;
        18: bitmap <= 590'b00100010001010010000010000100001001010100000101000001010000001101000010000010110100010010000011100100000100010101010100000000010101000100101010110010110101000101010101010001000110010100000001010101110000110101000001000100001000000000001010010100010000001001010011001011000000101010000001010101000100000100100100000000010100001100001010010000010101000110010000010001000010010000000011000000100000011100000010100000000001100000000001001000000000000001000010001110001000001100000001010010000000100000100000000000100111000000010000100000010100001001001001010001010110000000000010001000110001011;
        19: bitmap <= 590'b10011000000001010000010100100001000100000000101101000000000000010100100001011010000001010110000101010100000010100001000100000000100000000101101000010001001000000000000000010100010000010000000010000000000010110001001001000001001100000000011000010001000000001001000000001010000100010100000000100100000010100000000100000000100000000001010100000010000000010010010000000011010000000000000101000100010000010001010101100001000101000000001101010001000000001101010000010110000100010110000000110100000111010100000100000000000010000000111100010101001000000101000000011000010000010000000101001000000000;
        20: bitmap <= 590'b10001010000110001000011000100000010010000001010010001000100000010010100000010000100011000000000001001000000100101000100010000000101110000000100010001000101000000110100000000110001000001000000100011010001010000000100000100000101010100001001010000000100000000001001000101110100001001010000010100000000110101010000010000000101110100000101010001010011000000110001000010100001000001000000100100010001101001000000010000000010010000000100000000000100000010011000000010100100010100100000000000010000011000010100000000000101000100010100000000110101000000000100000001010001010000000000000100010001101;
        21: bitmap <= 590'b01010000011001010001000100000001010100000101000000000000000100000100000001000110100100010000000101010000010000000000000000010000010000000010010100000101010000010100000001000000000000000001000001000000010101010001000100000001010000000001000000000000000100000101000001100010000101010100000100010000010000000000000000010001000100000011010000010001010000000101000001000000000000000001000001010000010100101001010001000001000100000101000000000000010100000100000000110010100001010000000101010000010000000000000001010001000100000111010110010000010000010101000000000000000000000101000101010000010101;
        22: bitmap <= 590'b00101000001000111000100010100000001010000010000000000000000010001010100000100101100000101010000010000000001010000000000000100000001010000010011110001010000000000010100000101000000000000010100000101000001001011000101010100000100000000010000000000000001010001010000000001111100010100000000010001000000010000000000000101000101000000100101110001000000000000000000000101000000000000010000010101000011011110000101010000000100000000010100000000000001010000010100001001011000010001010000010001000001000000000000000101000100010000100001010001010001000000010100000001000000000000010100000001000001011;
        23: bitmap <= 590'b00000001010110001001010001010000000000010000000001010000000000000000000100011100100100010101000000000001010000000110010000010000000000010101010010000001010100000000000100000001001001000001000000000001000111001001010101010000000000010100000101010100000100000000000001001000000000010101000000000001010000010011010000000000000000010101100110010101010000000000000001000001011101000001000000000000000100011000000101010000000000010000000001110100000000000000000101001101100001010001000000000001000000010110010000010000000000010101110010000101000100000000000101000001011000000001000000000001000001;
        24: bitmap <= 590'b00000000101110011000101010001000000000001010000011001010000010000000000010101011100010100000100000000000001000001010101000001000000000001011001010001000101010000000000010100000111010100000100000000000100110110000001000001000000000001010000011100010000010000000000010101011100000101010100000000000101000001100101000001000000000000001100100001010101010000000000010100000101010100000100000000000100110000000001010101000000000001000000010001000000010000000000000110011000000001010100000000000101000000110001000001000000000000010101010001000101010000000000010000000011010100000100000000000101110;
        25: bitmap <= 590'b00000001010001000000000000000000101100000000010101111110000000000000000101010101000000000000000111111000000001011011001000000000000000010001000100000000000000011111100000000001101010100000000000000001010001010000000000000001111110000000010110111110000000000000000101000100000000000000000111111000000000010111010000000000000000010101010100000000000000011110100000000101110110100000000000000001010101010000000000000001111110000000010101110110000000000000000101000100000000000000000111101000000001011001111000000000000000000101010000000000000000011100100000000101111010100000000000000001010101;
        26: bitmap <= 590'b00000000001010101000000000000001111110000000001111111000000000000000000000101000000000000000000010110000000000101110111000000000000000001010101010000000000000001100100000000010111111100000000000000000101000101000000000000000110110000000000101111010000000000000000000101010100000000000000101101000000000111110111000000000000000001000101010000000000000011011100000000011101010100000000000000000101000101000000000000000110100000000001111111010000000000000000010101000100000000000000110111000000000011111100000000000000000001010101010000000000000010111100000000011001111100000000000000000101000;
        27: bitmap <= 590'b00010000010000000000000000010111101111010001010101011110000101000001000001000000000000000000011101111101000101010111101000010100000100000100000000000000000101111110110100010100011111100001010000010000010000000000000000010111111101010001010100111110000101000001000001000000000000000001011101111101000101010111011000010100000100000100000000000000000101011111110100010001011111100001010000010000010000000000000000010111111111010001010100111110000101000001000001000000000000000001011011101101000101010101111000010100000100000100000000000000000101111101110100010001011110000001010000010000010000;
        28: bitmap <= 590'b00001000001000000000000000000110111110101000101011111110000010100000100000100000000000000000111111101000100000101111111000001010000010000010000000000000000011111111101010001010110101100000101000001000001000000000000000001110111100101000101011011100000010100000100000100000000000000000101111110010100010101011111000001010000010000010000000000000000011111110101010001010111011100000101000001000001000000000000000001111111110001000101011111010000010100000100000100000000000000000101111111010100010101111101000001010000010000010000000000000000011011110101010001010111111100000101000001000001000;
        29: bitmap <= 590'b00010100000001010101010000010101111001000000000101010000000001000001010000000101010101000001010110110100000001010101000000010100000101000000010101010100000101001111010000000101010100000001010000010000000001010101010000010101111101000000010101010000000101000001010000000101010101000001010111010100000001010101000000010100000101000000010101010100000101011111010000000101010100000001000000010100000001010101010000010101111001000000010101000000000101000001010000000101010101000001010111110100000001010101000000000100000101000000010101010100000100011111010000000101010100000001010000010100000001;
        30: bitmap <= 590'b00001010000000101010101000001011111010100000001010101000000010100000101000000010101010100000101111101010000000101010100000001010000010100000001010101010000010111110101000000010101010000000101000001010000000101010101000001011111010100000001010101000000010100000101000000010101010100000101111101010000000101010100000001010000010100000001010101010000010110110101000000010101010000000101000000010000000101010101000001001111010100000001010101000000010100000101000000010101010100000101111100010000000101010100000001010000010100000001010101010000010111110101000000010101010000000101000001010000000;
        31: bitmap <= 590'b00010101000101010101000000000001010101000001000101010000000101010001010100010101010100000000000101010100000100000101000000010101000101010001010101010000000000010101010000010001010100000001010100010101000101010101000000000001010100000001000101010000000101010001010100010101010100000000000101010100000100010101000000010101000101010001010101010000000000010101010000010001010100000001010100010101000101010101000000000001010101000001000101010000000101010001010100010101010100000000000101010100000100010101000000010101000101010001010101010000000000010101010000010001010100000001010100010101000101;
        32: bitmap <= 590'b10001010100010101010100000000000101010100000100010101000000010101000101010001010101010000000000010101010000010001010100000001010100010101000101010101000000000001010101000001000101010000000101010001010100010101010100000000000101010100000100010101000000010101000101010001010101010000000000010101010000010001010100000001010100010101000101010101000000000001010101000001000101010000000101010001010100010101010100000000000101010100000100010101000000010101000101010001010101010000000000010101010000010001010100000001010100010101000101010101000000000001010101000001000101010000000101010001010100010;
        33: bitmap <= 590'b00010101000001010101000101000100010000000000010001010001000001010001010100000101010100010100010001000000000001000101000100000101000101010000010101010001010001000100000000000100010100010000010100010101000001010101000101000100010000000000010001010001000001010001010100000101010100010100010001000000000001000101000100000101000101010000010101010001010001000100000000000100010100010000010100010101000001010101000101000100010000000000010001010001000001010001010100000101010100010100010001000000000001000101000100000101000101010000010101010001010001000100000000000100010100010000010100010101000001;
        34: bitmap <= 590'b10001010100000101010100010100010001000000000001000101000100000101000101010000010101010001010001000100000000000100010100010000010100010101000001010101000101000100010000000000010001010001000001010001010100000101010100010100010001000000000001000101000100000101000101010000010101010001010001000100000000000100010100010000010100010101000001010101000101000100010000000000010001010001000001010001010100000101010100010100010001000000000001000101000100000101000101010000010101010001010001000100000000000100010100010000010100010101000001010101000101000100010000000000010001010001000001010001010100000;
        35: bitmap <= 590'b00000000000000000000000101000000000000011110000000000001010000000000000000000000000000010100000000000001111000000000000101000000000000000000000000000001010000000000000111100000000000010100000000000000000000000000000101000000000000011110000000000001010000000000000000000000000000010100000000000001111000000000000101000000000000000000000000000001010000000000000111100000000000010100000000000000000000000000000101000000000000011110000000000001010000000000000000000000000000010100000000000001111000000000000101000000000000000000000000000001010000000000000111100000000000010100000000000000000000;
        36: bitmap <= 590'b00000000000000000000000010100000000000011110000000000000101000000000000000000000000000001010000000000001111000000000000010100000000000000000000000000000101000000000000111100000000000001010000000000000000000000000000010100000000000011110000000000000101000000000000000000000000000001010000000000001111000000000000010100000000000000000000000000000101000000000000111100000000000001010000000000000000000000000000010100000000000011110000000000000101000000000000000000000000000001010000000000001111000000000000010100000000000000000000000000000101000000000000111100000000000001010000000000000000000;
        37: bitmap <= 590'b01011111000111110100000100000111110001010101000001010001010000010101111100011111010000010000011111000101010100000101000101000001010111110001111101000001000001111100010101010000010100010100000101011111000111110100000100000111110001010101000001010001010000010101111100011111010000010000011111000101010100000101000101000001010111110001111101000001000001111100010101010000010100010100000101011111000111110100000100000111110001010101000001010001010000010101111100011111010000010000011111000101010100000101000101000001010111110001111101000001000001111100010101010000010100010100000101011111000111;
        38: bitmap <= 590'b10111110100111101010000010000111101000101010100000101000101000001011111010011110101000001000011110100010101010000010100010100000101111101001111010100000100001111010001010101000001010001010000010111110100111101010000010000111101000101010100000101000101000001011111010011110101000001000011110100010101010000010100010100000101111101001111010100000100001111010001010101000001010001010000010111110100111101010000010000111101000101010100000101000101000001011111010011110101000001000011110100010101010000010100010100000101111101001111010100000100001111010001010101000001010001010000010111110100111;
        39: bitmap <= 590'b01010110000101111101000001010111110000010100000101010000000000000101011000010111110100000101011111000001010000010101000000000000010101100001011111010000010101111100000101000001010100000000000001010110000101111101000001010111110000010100000101010000000000000101011000010111110100000101011111000001010000010101000000000000010101100001011111010000010101111100000101000001010100000000000001010110000101111101000001010111110000010100000101010000000000000101011000010111110100000101011111000001010000010101000000000000010101100001011111010000010101111100000101000001010100000000000001010110000101;
        40: bitmap <= 590'b00101110000011111010100000101111101000001010000010101000000000000010111000001111101010000010111110100000101000001010100000000000001011100000111110101000001011111010000010100000101010000000000000101110000011111010100000101111101000001010000010101000000000000010111000001111101010000010111110100000101000001010100000000000001011100000111110101000001011111010000010100000101010000000000000101110000011111010100000101111101000001010000010101000000000000010111000001111101010000010111110100000101000001010100000000000001011100000111110101000001011111010000010100000101010000000000000101110000011;
        41: bitmap <= 590'b00010100000001000101000001000101010100000000000100000000000000000001010000000100010100000100010101010000000000010000000000000000000101000000010001010000010001010101000000000001000000000000000000010100000001000101000001000101010100000000000100000000000000000001010000000100010100000100010101010000000000010000000000000000000101000000010001010000010001010101000000000001000000000000000000010100000001000101000001000101010100000000000100000000000000000001010000000100010100000100010101010000000000010000000000000000000101000000010001010000010001010101000000000001000000000000000000010100000001;
        42: bitmap <= 590'b00001010000000100010100000100010101010000000000010000000000000000000101000000010001010000010001010101000000000001000000000000000000010100000001000101000001000101010100000000000100000000000000000001010000000100010100000100010101010000000000010000000000000000000101000000010001010000010001010101000000000001000000000000000000010100000001000101000001000101010100000000000100000000000000000001010000000100010100000100010101010000000000010000000000000000000101000000010001010000010001010101000000000001000000000000000000010100000001000101000001000101010100000000000100000000000000000001010000000;
        43: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        44: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        45: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        46: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        47: bitmap <= 590'b00000000000000000000101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        48: bitmap <= 590'b00000000000000000001111111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101;
        49: bitmap <= 590'b00000000000000000011111111101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        50: bitmap <= 590'b00000000000000000011111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        51: bitmap <= 590'b00000000000000000001111111101111111111111111111111111111111111111111111111111111111111111111111111111010101010101011101010101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010101010101110101010101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010101010111010101010101011111111111111111111111111111111111111111111111111111111111111111111;
        52: bitmap <= 590'b00000000000000000100011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        53: bitmap <= 590'b00000000000000000000001111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        54: bitmap <= 590'b00000000000000001000000111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        55: bitmap <= 590'b00000000000000001000001111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        56: bitmap <= 590'b00000000000000001000000111110111010000000000000000000000000000000000000000000000000000000000000111111111111111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111101111111111111111111000000000000000000000000000000000000000000000000000000000000000;
        57: bitmap <= 590'b00000000000000001000000011101111100000000000000000000000000000000000000000000000000000000000000010100000000000001110100000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000111010000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000011101000000000000011111000000000000000000000000000000000000000000000000000000000000000;
        58: bitmap <= 590'b00000000000000001000000111110111000000011111111111111111111111111111111000000000000000000000000111001111111111110110101111111111110111100000000000000000000000000111111111111111111111111111111111000001111111111111111111111111111111100001111111111111111111111111111111000000000000000000000000011100111111111111011010111111111111011110000000000000000000000000011111111111111111111111111111110000011111111111111111111111111111111000011111111111111111111111111111111100000000000000000000000001110011111111111101101011111111111101111000000000000000000000000001111111111111111111111111111111100000;
        59: bitmap <= 590'b00000000000000001000000011101111100000111111111111111111111111111111111000000000000000000000000010101111111111101110101111111111110111100000000000000000000000000111111111111111111111111111111110000011111111111111111111111111111111100001111111111111111111111111111111100000000000000000000000001010111111111110111010111111111111011110000000000000000000000000111111111111111111111111111111100000111111111111111111111111111111111000001111111111111111111111111111111100000000000000000000000000101011111111111011101011111111111101111000000000000000000000000001111111111111111111111111111111100000;
        60: bitmap <= 590'b00000000000000001000000111110111000000011111111111111111111111111111111000000000000000000000000111001111111111110110101111111111110111100000000000000000000000000111111111111111111111111111111111000001111111111111111111111111111111100001111111111111111111111111111111000000000000000000000000011100111111111111011010111111111111011110000000000000000000000000011111111111111111111111111111110000011111111111111111111111111111111000011111111111111111111111111111111100000000000000000000000001110011111111111101101011111111111101111000000000000000000000000001111111111111111111111111111111000000;
        61: bitmap <= 590'b00000000000000001000000011101111100000111111111111111111111111111111111000000000000000000000000010101111111111101110101111111111110111100000000000000000000000000111111111111111111111111111111110000011111111111111111111111111111111100001111111111111111111111111111111100000000000000000000000001010111111111110111010111111111111011110000000000000000000000000111111111111111111111111111111100000111111111111111111111111111111111000001111111111111111111111111111111100000000000000000000000000101011111111111011101011111111111101111000000000000000000000000001111111111111111111111111111111100000;
        62: bitmap <= 590'b00000000000000001000000111110111000000011111111111111111111111111111111000000000000000000000000111001111111111110110101111111111110111100000000000000000000000000111111111111111111111111111111111000001111111111111111111111111111111100001111111111111111111111111111111000000000000000000000000011100111111111111011010111111111111011110000000000000000000000000011111111111111111111111111111110000011111111111111111111111111111111000011111111111111111111111111111111100000000000000000000000001110011111111111101101011111111111101111000000000000000000000000001111111111111111111111111111111000000;
        63: bitmap <= 590'b00000000000000001000000011101111100000111111111111111111111111111111111000000000000000000000000010101111111111101110101111111111110111100000000000000000000000000111111111111111111111111111111110000011111111111111111111111111111111100001111111111111111111111111111111100000000000000000000000001010111111111110111010111111111111011110000000000000000000000000111111111111111111111111111111100000111111111111111111111111111111111000001111111111111111111111111111111100000000000000000000000000101011111111111011101011111111111101111000000000000000000000000001111111111111111111111111111111100000;
        64: bitmap <= 590'b00000000000000001000000111110111000000011111111111111111111111111111111000000000000000000000000111001111111111110110101111111111110111100000000000000000000000000111111111111111111111111111111111000001111111111111111111111111111111100001111111111111111111111111111111000000000000000000000000011100111111111111011010111111111111011110000000000000000000000000011111111111111111111111111111110000011111111111111111111111111111111000011111111111111111111111111111111100000000000000000000000001110011111111111101101011111111111101111000000000000000000000000001111111111111111111111111111111000000;
        65: bitmap <= 590'b00000000000000001000000011101111000000111111111111111111111111111111111000000000000000000000000010101111111111101110101111111111110111100000000000000000000000000111111111111111111111111111111110000011111111111111111111111111111111100001111111111111111111111111111111100000000000000000000000001010111111111110111010111111111111011110000000000000000000000000111111111111111111111111111111100000111111111111111111111111111111111000001111111111111111111111111111111100000000000000000000000000101011111111111011101011111111111101111000000000000000000000000001111111111111111111111111111111100000;
        66: bitmap <= 590'b00000000000000001000000111110111000000011111111111111111111111111111111000000000000000000000000111001111111111110110101111111111110111100000000000000000000000000111111111111111111111111111111111000001111111111111111111111111111111100001111111111111111111111111111111000000000000000000000000011100111111111111011010111111111111011110000000000000000000000000011111111111111111111111111111110000011111111111111111111111111111111000011111111111111111111111111111111100000000000000000000000001110011111111111101101011111111111101111000000000000000000000000001111111111111111111111111111111000000;
        67: bitmap <= 590'b00000000000000001000000011101111000000111111111111111111111111111111111000000000000000000000000010101111111111101110101111111111110111100000000000000000000000000111111111111111111111111111111110000011111111111111111111111111111111100001111111111111111111111111111111100000000000000000000000001010111111111110111010111111111111011110000000000000000000000000111111111111111111111111111111100000111111111111111111111111111111111000001111111111111111111111111111111100000000000000000000000000101011111111111011101011111111111101111000000000000000000000000001111111111111111111111111111111100000;
        68: bitmap <= 590'b00000000000000010000000111110111000000011111111111111111111111111111111000000000000000000000000111001111111111110110101111111111110111100000000000000000000000000111111111111111111111111111111111000001111111111111111111111111111111100001111111111111111111111111111111000000000000000000000000011100111111111111011010111111111111011110000000000000000000000000011111111111111111111111111111110000011111111111111111111111111111111000011111111111111111111111111111111100000000000000000000000001110011111111111101101011111111111101111000000000000000000000000001111111111111111111111111111111000000;
        69: bitmap <= 590'b00000000000000010000000011101111000000111111111111111111111111111111111000000000000000000000000010101111111111101110101111111111110111100000000000000000000000000111111111111111111111111111111110000011111111111111111111111111111111100001111111111111111111111111111111100000000000000000000000001010111111111110111010111111111111011110000000000000000000000000111111111111111111111111111111100000111111111111111111111111111111111000001111111111111111111111111111111100000000000000000000000000101011111111111011101011111111111101111000000000000000000000000001111111111111111111111111111111100000;
        70: bitmap <= 590'b00000000000000010000000111110111000000011111111111111111111111111111111000000000000000000000000111001111111111110110101111111111110111100000000000000000000000000111111111111111111111111111111111000001111111111111111111111111111111100001111111111111111111111111111111000000000000000000000000011100111111111111011010111111111111011110000000000000000000000000011111111111111111111111111111110000011111111111111111111111111111111000011111111111111111111111111111111100000000000000000000000001110011111111111101101011111111111101111000000000000000000000000001111111111111111111111111111111000000;
        71: bitmap <= 590'b00000000000000010000000011101111000000111111111111111111111111111111111000000000000000000000000010101111111111101110101111111111110111100000000000000000000000000111111111111111111111111111111110000011111111111111111111111111111111100001111111111111111111111111111111100000000000000000000000001010111111111110111010111111111111011110000000000000000000000000111111111111111111111111111111100000111111111111111111111111111111111000001111111111111111111111111111111100000000000000000000000000101011111111111011101011111111111101111000000000000000000000000001111111111111111111111111111111100000;
        72: bitmap <= 590'b00000000000000010000000111110111000000011111111111111111111111111111111000000000000000000000000111001111111111110110101111111111110111100000000000000000000000000111111111111111111111111111111111000001111111111111111111111111111111100001111111111111111111111111111111000000000000000000000000011100111111111111011010111111111111011110000000000000000000000000011111111111111111111111111111110000011111111111111111111111111111111000011111111111111111111111111111111100000000000000000000000001110011111111111101101011111111111101111000000000000000000000000001111111111111111111111111111111000000;
        73: bitmap <= 590'b00000000000000010000000011111111000000111111111111111111111111111111111000000000000000000000000010101111111111101110101111111111110111100000000000000000000000000111111111111111111111111111111110000011111111111111111111111111111111100001111111111111111111111111111111100000000000000000000000001010111111111110111010111111111111011110000000000000000000000000111111111111111111111111111111100000111111111111111111111111111111111000001111111111111111111111111111111100000000000000000000000000101011111111111011101011111111111101111000000000000000000000000001111111111111111111111111111111100000;
        74: bitmap <= 590'b00000000000000010000000111110111000000011111111111111111111111111111111000000000000000000000000111001111111111110110101111111111110111100000000000000000000000000111111111111111111111111111111111000001111111111111111111111111111111100001111111111111111111111111111111000000000000000000000000011100111111111111011010111111111111011110000000000000000000000000011111111111111111111111111111110000011111111111111111111111111111111000011111111111111111111111111111111100000000000000000000000001110011111111111101101011111111111101111000000000000000000000000001111111111111111111111111111111000000;
        75: bitmap <= 590'b00000000000000010000000011101111000000111111111111111111111111111111111000000000000000000000000010101111111111101110101111111111110111100000000000000000000000000111111111111111111111111111111110000011111111111111111111111111111111100001111111111111111111111111111111100000000000000000000000001010111111111110111010111111111111011110000000000000000000000000111111111111111111111111111111100000111111111111111111111111111111111000001111111111111111111111111111111100000000000000000000000000101011111111111011101011111111111101111000000000000000000000000001111111111111111111111111111111100000;
        76: bitmap <= 590'b00000000000000010000000111110111000000011111111111111111111111111111111000000000000000000000000111001111111111110110101111111111110111100000000000000000000000000111111111111111111111111111111111000001111111111111111111111111111111100001111111111111111111111111111111000000000000000000000000011100111111111111011010111111111111011110000000000000000000000000011111111111111111111111111111110000011111111111111111111111111111111000011111111111111111111111111111111100000000000000000000000001110011111111111101101011111111111101111000000000000000000000000001111111111111111111111111111111000000;
        77: bitmap <= 590'b00000000000000010000000011101111100000000000000000000000000000000000000000000000000000000000000010100000000000001110100000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000111010000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000011101000000000000011111000000000000000000000000000000000000000000000000000000000000000;
        78: bitmap <= 590'b00000000000000010000000111110111000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111111111111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111011111111111111110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111101111111111111111011000000000000000000000000000000000000000000000000000000000000000;
        79: bitmap <= 590'b00000000000000010000000011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111101111111111111111111111111111111111111111111111111111111111111111;
        80: bitmap <= 590'b00000000000000010000000111110111010101010101010101010101010101010101010101010101010101010101011111111111111111111100111111111111111101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111110011111111111111110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111111111111111111111001111111111111111010101010101010101010101010101010101010101010101010101010101010101;
        81: bitmap <= 590'b00000000000000010000000011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111101011111111111111111111111111111111111111111111111111111111111111;
        82: bitmap <= 590'b00000000000000010000000111110111010101010101010101010101010101010101010101010101010101010101011111111111111111111100111111111111111101011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111110011111111111111110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111111111111111111111001111111111111111010101010101010101010101010101010101010101010101010101010101010101;
        83: bitmap <= 590'b00000000000000010000000011101111101010101010101010101010101010101010101010101010101010101010101111111111111111111100111111111111111110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111111111111111111110011111111111111111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011111111111111111111001111111111111111101010101010101010101010101010101010101010101010101010101010101010;
        84: bitmap <= 590'b00000000000000010000000111110111010101010101010101010101010101010101010101010101010101010101011101111111111111111100111111111111111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111111111111111110011111111111111110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011111111111111111001111111111111111010101010101010101010101010101010101010101010101010101010101010101;
        85: bitmap <= 590'b00000000000000010000000011101111101010101010101010101010101010101010101010101010101010101010101111111111111111111100111111111111111110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111111111111111111110011111111111111111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011111111111111111111001111111111111111101010101010101010101010101010101010101010101010101010101010101010;
        86: bitmap <= 590'b00000000000000010000000111110111010101010101010101010101010101010101010101010101010101010101011101111111111111111100011111111111111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110111111111111111110001111111111111110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111011111111111111111000111111111111111010101010101010101010101010101010101010101010101010101010101010101;
        87: bitmap <= 590'b00000000000000010000001011101110101010101010101010101010101010101010101010101010101010101010101111111111111111111000111111111111111110111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111111111111111111100011111111111111111011101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011111111111111111110001111111111111111101110101010101010101010101010101010101010101010101010101010101010;
        88: bitmap <= 590'b00000000000000011000111111110111111101011101011101010101010101011101010101010101010101010111011101111111111111111100011111111111111101010101010101010101010101010101010101010101010101010101010101010101111111111101010101010101010111111101010101010101111111010101010111010101010101010101010101110111111111111111110001111111111111110101110101010101010101010101010101010101010101010101010101010101010101010101010101011101010101010101010101010101010101010101010101010101010101010101010101010111011111111111111111000111111111111111010111010101010101010101010101111101010101010101010101010111010111;
        89: bitmap <= 590'b00000000000000011111111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111101111111111111111111111111111111111111111111111111111111111111111;
        90: bitmap <= 590'b00000000000000010111000111110111111111111111111111111111111111111111111111111111111111111111111101111111111111111100011111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111110001111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111000111111111111111010111111111111111111111111111111111111111111111111111111111111111;
        91: bitmap <= 590'b00000000000000011000111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111101111111111111111111111111111111111111111111111111111111111111111;
        92: bitmap <= 590'b00000000000000010110111111110111010101010101010101010101010101010101010101010101010101010101011101011111111111111100011111111111111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110101111111111111110001111111111111110101110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010111111111111111000111111111111111010111010101010101010101010101010101010101010101010101010101010101;
        93: bitmap <= 590'b00000000000000011111111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111110101111111111111111111111111111111111111111111111111111111111111111;
        94: bitmap <= 590'b00000000000000010110111111111111010101010101010101010101010101010101010101010101010101010101011101011111111111111100010111111111111101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101110101111111111111110001011111111111110101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010111111111111111000101111111111111010101010101010101010101010101010101010101010101010101010101010101;
        95: bitmap <= 590'b00000000000000011111011011101110111111111111111111111111111111111111111111111111111111111111111111111010101010111000111010101010101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111101010101011100011101010101010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111110101010101110001110101010101010101111111111111111111111111111111111111111111111111111111111111111;
        96: bitmap <= 590'b00000000000000010111100111011101010101010101010101010101010101010101010101010101010101010101011101010101010101011100010101010101010101111101010101010101010101010101010101010101010101010101010101010101000101010101010001010101010101010101010101010101010101010101010101010101010101010001010101110101010101010101110001010101010101010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010001010101010111000101010101010111000101010101000101011101010100010001010101010101010101010101010101010101010101010101;
        97: bitmap <= 590'b00000000000000001000001011001110111101110111111111110111111111111011111011101111101111111011111111001010001010101000110010101010101010101111111011111111011111111111111111101110111111101111011110111111111110111011111111110110110111011110111011111110110111111011111011111011011110111111111010111010101010101010100011101010100010101011111111111111011111101111101111111111101111111101111011101111101111111101111011111011111110110111011111110111111111111101111011011111110111111111111101111010111010101010100010001110101000101010100110111011111111110111111111111111111111111111111111111111111111;
        98: bitmap <= 590'b00000000000000000011110111010101010101010101000100010101010001010101010101010101010101010101011001010101010100010000010101010101010111010100010101000101010101000100010101010101010001010101010101000101010101010101010101010101010101010101010101000101010101000101010100010101010101010100010101100101000100010100010000010101010100011101100100010001010101010101010100000101010001000101010101010101010100010101010101010100010101010101010001010101010100010101010101010100010100010100010101000111010101000100010101000100010101010101110111010101010101010100010001010101010101010101010101010101010101;
        99: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        100: bitmap <= 590'b10000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        101: bitmap <= 590'b00100101000110100100100101001000001001010101001010010000010000101010100100100100100001010000101010100001010101010101001000000100000100101001010010100101000001010100000001001001001001001000010101000010000101001000101010100100101001000010101010100101010010100100000101010100101010010010101001001001010101010010100001000001010010001001001010010101000001000010100100100010001001010000101001000010010100000101001000010010000100101001001000010000100101001001001010100010101010101010010100101001000010010010010000001001000101000001001001001010010010100100101000100001010000010100001000010010101001;
        102: bitmap <= 590'b00100010000010011001010100100101010101000000010000101010100101000000010100010010000001000101000000010100000000101000010010000010000001000110000100010000010110000100100100100100010100000101000000010100100010000100000000011010100100101001000000001000100000010011011000000010000001000100000010010110100010000100010010001000101000000000100001010010010010010000010101010010110010100011000101001001000011001000010100101101010001000010100101000101001000000001010010001100000100010000010010000101010000101000100100100100101010001000100100010010001000001001000000000000000101000001010001010000000010;
        103: bitmap <= 590'b10100001100001000100000010010000000000001000001100001000100000010001000101000101010000100100101100010101000100000110010001100001101000000001010100001010000010000010110000010010100001000100100010010010010001010001000100000001000000100000110001000100010100000001000100100010001001010010010001000000001001000001010100100100001010101010010000000001010001001010000000001000010000011000010000100101000000001000001010000000011000101000100101010000001001010100000001000000100010000101000001010000101000001010100010000010000000101010000001010001000010010001001101101010001000010101001100001010010001;
        104: bitmap <= 590'b00010100110000010000100000000110010100100101000010000000010101011000010000010001011000000010000101000001010010100000010100101000100011100000000100100001000011010000001001001000001010000100110001001010010100000100110001000000010100100100001001000001000110100001000010001001000101001000010000001001000100101000000010100000101010010010011010101000001100101000100101000010010010000000000100010001101101001001000001000000000010100100000100001001000101000010010000010101010001100100010100001000101010000000101010001000100101000101010100000101010010001000100000101001000010000000000101000001001000;
        105: bitmap <= 590'b00000000001001000010010101010000000001000010010001001100100000000010000101000000000000100100100000000100000000000001000000000010000100001010000010000100101000001010001100000001001001010001001000100001000001010010000100011000100000001000100100010000000001001000010100010000100000100101001010010010000000000010010000010101000000000000000001000010010000000001000000001000000010010101001001000000000000100010001000010101010000000000100000000100010000010000101010100100000000010000100001000100000001011000000000100000010000010000101001000000001000010010001010000000001001101000100000001000100010;
        106: bitmap <= 590'b11010010100100001001000000001000101010100000001000100010010100000000000000101000010001010000001001001010010010001010000101001000001000000001001000000000000000100000100000101000100100000000000100000100001000001001000001000000010010100100001000001001010000000100000010000100010000000000100001000000010001001001000100000000000101000010100000100000100001000100001100100010010000000000010000101010001010001000100100100010000010000010010100100010000100000100000000000001010000000010000100100000100100000100101010101001000010000000000000101010000001001000100000001011000100000010001000100110000100;
        107: bitmap <= 590'b00000000000010000000100000000000000000010000000000000000000010010100100000001010000000000010000000100001000000000000100000000100100001000000010001100010010000000000000000000000000010000100000100000010000010000000000000000100001000000010000100101000001000100010000000100000010010100000000000001010010001000000100010010101000000010000000000100000000000100000100000010000000000010100001000000000000000000000000000100000001001000000000000100000000000000010000100100000010000000000010000000100000000000000000000001000000000010000000000000001000000000000010000000000100000000000001000000001000000;
        108: bitmap <= 590'b01000000000000000000000100001000000001000100000000000000010000000010000100000000101000010000000000000000000100100000000000000000000000101000000000000000001000100010000000000000000001000001000000000000000000000010100010000000000000000000000000000000100000000010000100000000000000000000010000000000000000000000000000000000000000000001010000010000001000001000000000000100010100000000000000000000000000001000000000000010000000010000000000001001000100000001000000000000000100010000000000010000000000000001000000000000100000001000000000000000000000000000001000000000000010010000000001000000000010;
        109: bitmap <= 590'b00001001000000000000000001000100000100000000010000101000000000000000000000000000000000000000100000000000010000000000000000000010000000000001000000001000000000000100000100010000000000000000000000010000000000100000000000000000000010000000000010000000000100000000000000010000100000000100001001000000000000000100000000000000000100010000000000000010000000000000001000010000000000000001000000000100100000100000100000001000000000100000010100000000000000100000000000000000100000000010000001000000010010000100000000000010000010000000010000000100100100000100000000000000000000000001000100000000000000;
        110: bitmap <= 590'b00000000000010101000000000000000000000000001000000000000000100000000100000000000000100000000010000000000000000010000010001000000010000000000000001000000000000000000000000000010000000000000001000000000000000000000010000000100000000000000100000000010000000000000010000000100000001000000000000000001000000100000001000000001000000000000000000000000000000000000000000000000000000000000000010000000000100000000000001000000000000000001000000000000100000000000001000000000000001000000001000000000001000000000000100001000001000000010001000100000000001000000000000010100000000001000000000000000001000;
        111: bitmap <= 590'b00000000000000000010000000000000000000000000000000000000000010000000000000000000000000010000000001000000000000000000010000000000000000000000000000000001000000000001000000000000000010000000000000001000010000000000001000000100000000000000000000000000000010000100000000000000000000000100000000000000000000000000000100000000000000001000000000000000000000000010000000000000000001000000000000000000000000000000000000000000001000000000000000000000000100000000000000100000100000000000000000000000000000000000000010000000000000100000000000000000000000100000000010000010000000000000000000010000000000;
        112: bitmap <= 590'b00000000100000000000000000000000000000100000100000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000;
        113: bitmap <= 590'b00000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        114: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000010000000000100000000000000000010000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        115: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        116: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        117: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        118: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        119: bitmap <= 590'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

    default: bitmap <= 0;
       endcase
 end
        endmodule