module bannerword4_12 (
    input wire clk,  // clock
    input wire [4:0] address,  // reset
    output reg [70:0] outdata
  );
  
  (* rom_style = "block" *)
  
  reg [4:0] address_reg;

  /* Combinational Logic */
  always @* begin
    case(address_reg)
      0: outdata = 71'b00000000000000000111111000111111111000111111000000111111000000111111111;
      1: outdata = 71'b00000000000000000111111000111111111000111111000000111111000000111111111;
      2: outdata = 71'b00000000000000000111111000111111111000111111000000111111000000111111111;
      3: outdata = 71'b11000000000000111000000000000111000000111000111000111000111000000111000;
      4: outdata = 71'b11000000000000111000000000000111000000111000111000111000111000000111000;
      5: outdata = 71'b11000000000000111000000000000111000000111000111000111000111000000111000;
      6: outdata = 71'b11000000000000000111000000000111000000111111111000111111000000000111000;
      7: outdata = 71'b11000000000000000111000000000111000000111111111000111111000000000111000;
      8: outdata = 71'b11000000000000000111000000000111000000111111111000111111000000000111000;
      9: outdata = 71'b11000000000000000000111000000111000000111000111000111000111000000111000;
      10: outdata = 71'b11000000000000000000111000000111000000111000111000111000111000000111000;
      11: outdata = 71'b11000000000000000000111000000111000000111000111000111000111000000111000;
      12: outdata = 71'b11000000000000111111111000000111000000111000111000111000111000000111000;
      13: outdata = 71'b11000000000000111111111000000111000000111000111000111000111000000111000;
      14: outdata = 71'b11000000000000111111111000000111000000111000111000111000111000000111000;
    default: outdata = 0;
    endcase
  end
  
  /* Sequential Logic */
  always @(posedge clk) begin
    address_reg <= address;
  end
  
endmodule